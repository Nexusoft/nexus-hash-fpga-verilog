// Created by cells_xtra.py from Xilinx models

module FDCE (...);
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] INIT = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_CLR_INVERTED" *)
    input CLR;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
endmodule

module FDPE (...);
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] IS_PRE_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    (* invertible_pin = "IS_PRE_INVERTED" *)
    input PRE;
endmodule

module FDRE (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] IS_R_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    (* invertible_pin = "IS_R_INVERTED" *)
    input R;
endmodule

module FDSE (...);
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] IS_S_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    (* invertible_pin = "IS_S_INVERTED" *)
    input S;
endmodule

module LDCE (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    (* invertible_pin = "IS_CLR_INVERTED" *)
    input CLR;
    input D;
    (* invertible_pin = "IS_G_INVERTED" *)
    input G;
    input GE;
endmodule

module LDPE (...);
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_G_INVERTED = 1'b0;
    parameter [0:0] IS_PRE_INVERTED = 1'b0;
    parameter MSGON = "TRUE";
    parameter XON = "TRUE";
    output Q;
    input D;
    (* invertible_pin = "IS_G_INVERTED" *)
    input G;
    input GE;
    (* invertible_pin = "IS_PRE_INVERTED" *)
    input PRE;
endmodule

module AND2B1L (...);
    parameter [0:0] IS_SRI_INVERTED = 1'b0;
    output O;
    input DI;
    (* invertible_pin = "IS_SRI_INVERTED" *)
    input SRI;
endmodule

module OR2L (...);
    parameter [0:0] IS_SRI_INVERTED = 1'b0;
    output O;
    input DI;
    (* invertible_pin = "IS_SRI_INVERTED" *)
    input SRI;
endmodule

module LUT1 (...);
    parameter [1:0] INIT = 2'h0;
    input I0;
    output O;
endmodule

module LUT2 (...);
    parameter [3:0] INIT = 4'h0;
    input I0;
    input I1;
    output O;
endmodule

module LUT3 (...);
    parameter [7:0] INIT = 8'h00;
    input I0;
    input I1;
    input I2;
    output O;
endmodule

module LUT4 (...);
    parameter [15:0] INIT = 16'h0000;
    input I0;
    input I1;
    input I2;
    input I3;
    output O;
endmodule

module LUT5 (...);
    parameter [31:0] INIT = 32'h00000000;
    input I0;
    input I1;
    input I2;
    input I3;
    input I4;
    output O;
endmodule

module LUT6 (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    input I0;
    input I1;
    input I2;
    input I3;
    input I4;
    input I5;
    output O;
endmodule

module LUT6_2 (...);
    parameter [63:0] INIT = 64'h0000000000000000;
    input I0;
    input I1;
    input I2;
    input I3;
    input I4;
    input I5;
    output O5;
    output O6;
endmodule

module MUXF5 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module MUXF6 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module MUXF7 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module MUXF8 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module MUXF9 (...);
    output O;
    input I0;
    input I1;
    input S;
endmodule

module CARRY4 (...);
    output [3:0] CO;
    output [3:0] O;
    input CI;
    input CYINIT;
    input [3:0] DI;
    input [3:0] S;
endmodule

module CARRY8 (...);
    parameter CARRY_TYPE = "SINGLE_CY8";
    output [7:0] CO;
    output [7:0] O;
    input CI;
    input CI_TOP;
    input [7:0] DI;
    input [7:0] S;
endmodule

module MUXCY (...);
    output O;
    input CI;
    input DI;
    input S;
endmodule

module XORCY (...);
    output O;
    input CI;
    input LI;
endmodule

module SRL16 (...);
    parameter [15:0] INIT = 16'h0000;
    output Q;
    input A0;
    input A1;
    input A2;
    input A3;
    (* clkbuf_sink *)
    input CLK;
    input D;
endmodule

module SRL16E (...);
    parameter [15:0] INIT = 16'h0000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output Q;
    input A0;
    input A1;
    input A2;
    input A3;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input D;
endmodule

module SRLC16 (...);
    parameter [15:0] INIT = 16'h0000;
    output Q;
    output Q15;
    input A0;
    input A1;
    input A2;
    input A3;
    (* clkbuf_sink *)
    input CLK;
    input D;
endmodule

module SRLC16E (...);
    parameter [15:0] INIT = 16'h0000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output Q;
    output Q15;
    input A0;
    input A1;
    input A2;
    input A3;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input D;
endmodule

module SRLC32E (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output Q;
    output Q31;
    input [4:0] A;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input D;
endmodule

module CFGLUT5 (...);
    parameter [31:0] INIT = 32'h00000000;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    output CDO;
    output O5;
    output O6;
    input I4;
    input I3;
    input I2;
    input I1;
    input I0;
    input CDI;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
endmodule

module FIFO18E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO18";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 36'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 36'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output [31:0] DO;
    output [3:0] DOP;
    output EMPTY;
    output FULL;
    output [11:0] RDCOUNT;
    output RDERR;
    output [11:0] WRCOUNT;
    output WRERR;
    input [31:0] DI;
    input [3:0] DIP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO36E1 (...);
    parameter ALMOST_EMPTY_OFFSET = 13'h0080;
    parameter ALMOST_FULL_OFFSET = 13'h0080;
    parameter integer DATA_WIDTH = 4;
    parameter integer DO_REG = 1;
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter EN_SYN = "FALSE";
    parameter FIFO_MODE = "FIFO36";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter INIT = 72'h0;
    parameter SIM_DEVICE = "VIRTEX6";
    parameter SRVAL = 72'h0;
    parameter IS_RDCLK_INVERTED = 1'b0;
    parameter IS_RDEN_INVERTED = 1'b0;
    parameter IS_RSTREG_INVERTED = 1'b0;
    parameter IS_RST_INVERTED = 1'b0;
    parameter IS_WRCLK_INVERTED = 1'b0;
    parameter IS_WREN_INVERTED = 1'b0;
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output DBITERR;
    output [63:0] DO;
    output [7:0] DOP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output SBITERR;
    output [12:0] WRCOUNT;
    output WRERR;
    input [63:0] DI;
    input [7:0] DIP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO18E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [35:0] INIT = 36'h000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL = 36'h000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [31:0] CASDOUT;
    output [3:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output [31:0] DOUT;
    output [3:0] DOUTP;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [12:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output [12:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [31:0] CASDIN;
    input [3:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [31:0] DIN;
    input [3:0] DINP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module FIFO36E2 (...);
    parameter CASCADE_ORDER = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter FIRST_WORD_FALL_THROUGH = "FALSE";
    parameter [71:0] INIT = 72'h000000000000000000;
    parameter [0:0] IS_RDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RDEN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_WRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_WREN_INVERTED = 1'b0;
    parameter integer PROG_EMPTY_THRESH = 256;
    parameter integer PROG_FULL_THRESH = 256;
    parameter RDCOUNT_TYPE = "RAW_PNTR";
    parameter integer READ_WIDTH = 4;
    parameter REGISTER_MODE = "UNREGISTERED";
    parameter RSTREG_PRIORITY = "RSTREG";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [71:0] SRVAL = 72'h000000000000000000;
    parameter WRCOUNT_TYPE = "RAW_PNTR";
    parameter integer WRITE_WIDTH = 4;
    output [63:0] CASDOUT;
    output [7:0] CASDOUTP;
    output CASNXTEMPTY;
    output CASPRVRDEN;
    output DBITERR;
    output [63:0] DOUT;
    output [7:0] DOUTP;
    output [7:0] ECCPARITY;
    output EMPTY;
    output FULL;
    output PROGEMPTY;
    output PROGFULL;
    output [13:0] RDCOUNT;
    output RDERR;
    output RDRSTBUSY;
    output SBITERR;
    output [13:0] WRCOUNT;
    output WRERR;
    output WRRSTBUSY;
    input [63:0] CASDIN;
    input [7:0] CASDINP;
    input CASDOMUX;
    input CASDOMUXEN;
    input CASNXTRDEN;
    input CASOREGIMUX;
    input CASOREGIMUXEN;
    input CASPRVEMPTY;
    input [63:0] DIN;
    input [7:0] DINP;
    input INJECTDBITERR;
    input INJECTSBITERR;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_RDCLK_INVERTED" *)
    input RDCLK;
    (* invertible_pin = "IS_RDEN_INVERTED" *)
    input RDEN;
    input REGCE;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RSTREG_INVERTED" *)
    input RSTREG;
    input SLEEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_WRCLK_INVERTED" *)
    input WRCLK;
    (* invertible_pin = "IS_WREN_INVERTED" *)
    input WREN;
endmodule

module RAMB18E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [17:0] INIT_A = 18'h00000;
    parameter [17:0] INIT_B = 18'h00000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [17:0] SRVAL_A = 18'h00000;
    parameter [17:0] SRVAL_B = 18'h00000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [15:0] CASDOUTA;
    output [15:0] CASDOUTB;
    output [1:0] CASDOUTPA;
    output [1:0] CASDOUTPB;
    output [15:0] DOUTADOUT;
    output [15:0] DOUTBDOUT;
    output [1:0] DOUTPADOUTP;
    output [1:0] DOUTPBDOUTP;
    input [13:0] ADDRARDADDR;
    input [13:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [15:0] CASDINA;
    input [15:0] CASDINB;
    input [1:0] CASDINPA;
    input [1:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKARDCLK_INVERTED" *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKBWRCLK_INVERTED" *)
    input CLKBWRCLK;
    input [15:0] DINADIN;
    input [15:0] DINBDIN;
    input [1:0] DINPADINP;
    input [1:0] DINPBDINP;
    (* invertible_pin = "IS_ENARDEN_INVERTED" *)
    input ENARDEN;
    (* invertible_pin = "IS_ENBWREN_INVERTED" *)
    input ENBWREN;
    input REGCEAREGCE;
    input REGCEB;
    (* invertible_pin = "IS_RSTRAMARSTRAM_INVERTED" *)
    input RSTRAMARSTRAM;
    (* invertible_pin = "IS_RSTRAMB_INVERTED" *)
    input RSTRAMB;
    (* invertible_pin = "IS_RSTREGARSTREG_INVERTED" *)
    input RSTREGARSTREG;
    (* invertible_pin = "IS_RSTREGB_INVERTED" *)
    input RSTREGB;
    input SLEEP;
    input [1:0] WEA;
    input [3:0] WEBWE;
endmodule

module RAMB36E2 (...);
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter CLOCK_DOMAINS = "INDEPENDENT";
    parameter integer DOA_REG = 1;
    parameter integer DOB_REG = 1;
    parameter ENADDRENA = "FALSE";
    parameter ENADDRENB = "FALSE";
    parameter EN_ECC_PIPE = "FALSE";
    parameter EN_ECC_READ = "FALSE";
    parameter EN_ECC_WRITE = "FALSE";
    parameter [255:0] INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INITP_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_40 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_41 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_42 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_43 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_44 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_45 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_46 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_47 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_48 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_49 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_4F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_50 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_51 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_52 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_53 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_54 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_55 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_56 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_57 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_58 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_59 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_5F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_60 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_61 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_62 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_63 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_64 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_65 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_66 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_67 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_68 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_69 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_6F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_70 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_71 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_72 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_73 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_74 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_75 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_76 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_77 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_78 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_79 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [255:0] INIT_7F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter [35:0] INIT_A = 36'h000000000;
    parameter [35:0] INIT_B = 36'h000000000;
    parameter INIT_FILE = "NONE";
    parameter [0:0] IS_CLKARDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_CLKBWRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_ENARDEN_INVERTED = 1'b0;
    parameter [0:0] IS_ENBWREN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMARSTRAM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTRAMB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGARSTREG_INVERTED = 1'b0;
    parameter [0:0] IS_RSTREGB_INVERTED = 1'b0;
    parameter RDADDRCHANGEA = "FALSE";
    parameter RDADDRCHANGEB = "FALSE";
    parameter integer READ_WIDTH_A = 0;
    parameter integer READ_WIDTH_B = 0;
    parameter RSTREG_PRIORITY_A = "RSTREG";
    parameter RSTREG_PRIORITY_B = "RSTREG";
    parameter SIM_COLLISION_CHECK = "ALL";
    parameter SLEEP_ASYNC = "FALSE";
    parameter [35:0] SRVAL_A = 36'h000000000;
    parameter [35:0] SRVAL_B = 36'h000000000;
    parameter WRITE_MODE_A = "NO_CHANGE";
    parameter WRITE_MODE_B = "NO_CHANGE";
    parameter integer WRITE_WIDTH_A = 0;
    parameter integer WRITE_WIDTH_B = 0;
    output [31:0] CASDOUTA;
    output [31:0] CASDOUTB;
    output [3:0] CASDOUTPA;
    output [3:0] CASDOUTPB;
    output CASOUTDBITERR;
    output CASOUTSBITERR;
    output DBITERR;
    output [31:0] DOUTADOUT;
    output [31:0] DOUTBDOUT;
    output [3:0] DOUTPADOUTP;
    output [3:0] DOUTPBDOUTP;
    output [7:0] ECCPARITY;
    output [8:0] RDADDRECC;
    output SBITERR;
    input [14:0] ADDRARDADDR;
    input [14:0] ADDRBWRADDR;
    input ADDRENA;
    input ADDRENB;
    input CASDIMUXA;
    input CASDIMUXB;
    input [31:0] CASDINA;
    input [31:0] CASDINB;
    input [3:0] CASDINPA;
    input [3:0] CASDINPB;
    input CASDOMUXA;
    input CASDOMUXB;
    input CASDOMUXEN_A;
    input CASDOMUXEN_B;
    input CASINDBITERR;
    input CASINSBITERR;
    input CASOREGIMUXA;
    input CASOREGIMUXB;
    input CASOREGIMUXEN_A;
    input CASOREGIMUXEN_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKARDCLK_INVERTED" *)
    input CLKARDCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKBWRCLK_INVERTED" *)
    input CLKBWRCLK;
    input [31:0] DINADIN;
    input [31:0] DINBDIN;
    input [3:0] DINPADINP;
    input [3:0] DINPBDINP;
    input ECCPIPECE;
    (* invertible_pin = "IS_ENARDEN_INVERTED" *)
    input ENARDEN;
    (* invertible_pin = "IS_ENBWREN_INVERTED" *)
    input ENBWREN;
    input INJECTDBITERR;
    input INJECTSBITERR;
    input REGCEAREGCE;
    input REGCEB;
    (* invertible_pin = "IS_RSTRAMARSTRAM_INVERTED" *)
    input RSTRAMARSTRAM;
    (* invertible_pin = "IS_RSTRAMB_INVERTED" *)
    input RSTRAMB;
    (* invertible_pin = "IS_RSTREGARSTREG_INVERTED" *)
    input RSTREGARSTREG;
    (* invertible_pin = "IS_RSTREGB_INVERTED" *)
    input RSTREGB;
    input SLEEP;
    input [3:0] WEA;
    input [7:0] WEBWE;
endmodule

module URAM288 (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter CASCADE_ORDER_A = "NONE";
    parameter CASCADE_ORDER_B = "NONE";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter MATRIX_ID = "NONE";
    parameter integer NUM_UNIQUE_SELF_ADDR_A = 1;
    parameter integer NUM_UNIQUE_SELF_ADDR_B = 1;
    parameter integer NUM_URAM_IN_MATRIX = 1;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter REG_CAS_A = "FALSE";
    parameter REG_CAS_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter [10:0] SELF_ADDR_A = 11'h000;
    parameter [10:0] SELF_ADDR_B = 11'h000;
    parameter [10:0] SELF_MASK_A = 11'h7FF;
    parameter [10:0] SELF_MASK_B = 11'h7FF;
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output [22:0] CAS_OUT_ADDR_A;
    output [22:0] CAS_OUT_ADDR_B;
    output [8:0] CAS_OUT_BWE_A;
    output [8:0] CAS_OUT_BWE_B;
    output CAS_OUT_DBITERR_A;
    output CAS_OUT_DBITERR_B;
    output [71:0] CAS_OUT_DIN_A;
    output [71:0] CAS_OUT_DIN_B;
    output [71:0] CAS_OUT_DOUT_A;
    output [71:0] CAS_OUT_DOUT_B;
    output CAS_OUT_EN_A;
    output CAS_OUT_EN_B;
    output CAS_OUT_RDACCESS_A;
    output CAS_OUT_RDACCESS_B;
    output CAS_OUT_RDB_WR_A;
    output CAS_OUT_RDB_WR_B;
    output CAS_OUT_SBITERR_A;
    output CAS_OUT_SBITERR_B;
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output RDACCESS_A;
    output RDACCESS_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    input [22:0] CAS_IN_ADDR_A;
    input [22:0] CAS_IN_ADDR_B;
    input [8:0] CAS_IN_BWE_A;
    input [8:0] CAS_IN_BWE_B;
    input CAS_IN_DBITERR_A;
    input CAS_IN_DBITERR_B;
    input [71:0] CAS_IN_DIN_A;
    input [71:0] CAS_IN_DIN_B;
    input [71:0] CAS_IN_DOUT_A;
    input [71:0] CAS_IN_DOUT_B;
    input CAS_IN_EN_A;
    input CAS_IN_EN_B;
    input CAS_IN_RDACCESS_A;
    input CAS_IN_RDACCESS_B;
    input CAS_IN_RDB_WR_A;
    input CAS_IN_RDB_WR_B;
    input CAS_IN_SBITERR_A;
    input CAS_IN_SBITERR_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    (* invertible_pin = "IS_EN_A_INVERTED" *)
    input EN_A;
    (* invertible_pin = "IS_EN_B_INVERTED" *)
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    (* invertible_pin = "IS_RDB_WR_A_INVERTED" *)
    input RDB_WR_A;
    (* invertible_pin = "IS_RDB_WR_B_INVERTED" *)
    input RDB_WR_B;
    (* invertible_pin = "IS_RST_A_INVERTED" *)
    input RST_A;
    (* invertible_pin = "IS_RST_B_INVERTED" *)
    input RST_B;
    input SLEEP;
endmodule

module URAM288_BASE (...);
    parameter integer AUTO_SLEEP_LATENCY = 8;
    parameter integer AVG_CONS_INACTIVE_CYCLES = 10;
    parameter BWE_MODE_A = "PARITY_INTERLEAVED";
    parameter BWE_MODE_B = "PARITY_INTERLEAVED";
    parameter EN_AUTO_SLEEP_MODE = "FALSE";
    parameter EN_ECC_RD_A = "FALSE";
    parameter EN_ECC_RD_B = "FALSE";
    parameter EN_ECC_WR_A = "FALSE";
    parameter EN_ECC_WR_B = "FALSE";
    parameter IREG_PRE_A = "FALSE";
    parameter IREG_PRE_B = "FALSE";
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_EN_A_INVERTED = 1'b0;
    parameter [0:0] IS_EN_B_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_A_INVERTED = 1'b0;
    parameter [0:0] IS_RDB_WR_B_INVERTED = 1'b0;
    parameter [0:0] IS_RST_A_INVERTED = 1'b0;
    parameter [0:0] IS_RST_B_INVERTED = 1'b0;
    parameter OREG_A = "FALSE";
    parameter OREG_B = "FALSE";
    parameter OREG_ECC_A = "FALSE";
    parameter OREG_ECC_B = "FALSE";
    parameter RST_MODE_A = "SYNC";
    parameter RST_MODE_B = "SYNC";
    parameter USE_EXT_CE_A = "FALSE";
    parameter USE_EXT_CE_B = "FALSE";
    output DBITERR_A;
    output DBITERR_B;
    output [71:0] DOUT_A;
    output [71:0] DOUT_B;
    output SBITERR_A;
    output SBITERR_B;
    input [22:0] ADDR_A;
    input [22:0] ADDR_B;
    input [8:0] BWE_A;
    input [8:0] BWE_B;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [71:0] DIN_A;
    input [71:0] DIN_B;
    (* invertible_pin = "IS_EN_A_INVERTED" *)
    input EN_A;
    (* invertible_pin = "IS_EN_B_INVERTED" *)
    input EN_B;
    input INJECT_DBITERR_A;
    input INJECT_DBITERR_B;
    input INJECT_SBITERR_A;
    input INJECT_SBITERR_B;
    input OREG_CE_A;
    input OREG_CE_B;
    input OREG_ECC_CE_A;
    input OREG_ECC_CE_B;
    (* invertible_pin = "IS_RDB_WR_A_INVERTED" *)
    input RDB_WR_A;
    (* invertible_pin = "IS_RDB_WR_B_INVERTED" *)
    input RDB_WR_B;
    (* invertible_pin = "IS_RST_A_INVERTED" *)
    input RST_A;
    (* invertible_pin = "IS_RST_B_INVERTED" *)
    input RST_B;
    input SLEEP;
endmodule

module DSP48E1 (...);
    parameter integer ACASCREG = 1;
    parameter integer ADREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter integer AREG = 1;
    parameter AUTORESET_PATDET = "NO_RESET";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter integer DREG = 1;
    parameter integer INMODEREG = 1;
    parameter integer MREG = 1;
    parameter integer OPMODEREG = 1;
    parameter integer PREG = 1;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter USE_DPORT = "FALSE";
    parameter USE_MULT = "MULTIPLY";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter [3:0] IS_ALUMODE_INVERTED = 4'b0;
    parameter [0:0] IS_CARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [4:0] IS_INMODE_INVERTED = 5'b0;
    parameter [6:0] IS_OPMODE_INVERTED = 7'b0;
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    input [29:0] A;
    input [29:0] ACIN;
    (* invertible_pin = "IS_ALUMODE_INVERTED" *)
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    (* invertible_pin = "IS_CARRYIN_INVERTED" *)
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEAD;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CED;
    input CEINMODE;
    input CEM;
    input CEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [24:0] D;
    (* invertible_pin = "IS_INMODE_INVERTED" *)
    input [4:0] INMODE;
    input MULTSIGNIN;
    (* invertible_pin = "IS_OPMODE_INVERTED" *)
    input [6:0] OPMODE;
    input [47:0] PCIN;
    input RSTA;
    input RSTALLCARRYIN;
    input RSTALUMODE;
    input RSTB;
    input RSTC;
    input RSTCTRL;
    input RSTD;
    input RSTINMODE;
    input RSTM;
    input RSTP;
endmodule

module DSP48E2 (...);
    parameter integer ACASCREG = 1;
    parameter integer ADREG = 1;
    parameter integer ALUMODEREG = 1;
    parameter AMULTSEL = "A";
    parameter integer AREG = 1;
    parameter AUTORESET_PATDET = "NO_RESET";
    parameter AUTORESET_PRIORITY = "RESET";
    parameter A_INPUT = "DIRECT";
    parameter integer BCASCREG = 1;
    parameter BMULTSEL = "B";
    parameter integer BREG = 1;
    parameter B_INPUT = "DIRECT";
    parameter integer CARRYINREG = 1;
    parameter integer CARRYINSELREG = 1;
    parameter integer CREG = 1;
    parameter integer DREG = 1;
    parameter integer INMODEREG = 1;
    parameter [3:0] IS_ALUMODE_INVERTED = 4'b0000;
    parameter [0:0] IS_CARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [4:0] IS_INMODE_INVERTED = 5'b00000;
    parameter [8:0] IS_OPMODE_INVERTED = 9'b000000000;
    parameter [0:0] IS_RSTALLCARRYIN_INVERTED = 1'b0;
    parameter [0:0] IS_RSTALUMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTA_INVERTED = 1'b0;
    parameter [0:0] IS_RSTB_INVERTED = 1'b0;
    parameter [0:0] IS_RSTCTRL_INVERTED = 1'b0;
    parameter [0:0] IS_RSTC_INVERTED = 1'b0;
    parameter [0:0] IS_RSTD_INVERTED = 1'b0;
    parameter [0:0] IS_RSTINMODE_INVERTED = 1'b0;
    parameter [0:0] IS_RSTM_INVERTED = 1'b0;
    parameter [0:0] IS_RSTP_INVERTED = 1'b0;
    parameter [47:0] MASK = 48'h3FFFFFFFFFFF;
    parameter integer MREG = 1;
    parameter integer OPMODEREG = 1;
    parameter [47:0] PATTERN = 48'h000000000000;
    parameter PREADDINSEL = "A";
    parameter integer PREG = 1;
    parameter [47:0] RND = 48'h000000000000;
    parameter SEL_MASK = "MASK";
    parameter SEL_PATTERN = "PATTERN";
    parameter USE_MULT = "MULTIPLY";
    parameter USE_PATTERN_DETECT = "NO_PATDET";
    parameter USE_SIMD = "ONE48";
    parameter USE_WIDEXOR = "FALSE";
    parameter XORSIMD = "XOR24_48_96";
    output [29:0] ACOUT;
    output [17:0] BCOUT;
    output CARRYCASCOUT;
    output [3:0] CARRYOUT;
    output MULTSIGNOUT;
    output OVERFLOW;
    output [47:0] P;
    output PATTERNBDETECT;
    output PATTERNDETECT;
    output [47:0] PCOUT;
    output UNDERFLOW;
    output [7:0] XOROUT;
    input [29:0] A;
    input [29:0] ACIN;
    (* invertible_pin = "IS_ALUMODE_INVERTED" *)
    input [3:0] ALUMODE;
    input [17:0] B;
    input [17:0] BCIN;
    input [47:0] C;
    input CARRYCASCIN;
    (* invertible_pin = "IS_CARRYIN_INVERTED" *)
    input CARRYIN;
    input [2:0] CARRYINSEL;
    input CEA1;
    input CEA2;
    input CEAD;
    input CEALUMODE;
    input CEB1;
    input CEB2;
    input CEC;
    input CECARRYIN;
    input CECTRL;
    input CED;
    input CEINMODE;
    input CEM;
    input CEP;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [26:0] D;
    (* invertible_pin = "IS_INMODE_INVERTED" *)
    input [4:0] INMODE;
    input MULTSIGNIN;
    (* invertible_pin = "IS_OPMODE_INVERTED" *)
    input [8:0] OPMODE;
    input [47:0] PCIN;
    (* invertible_pin = "IS_RSTA_INVERTED" *)
    input RSTA;
    (* invertible_pin = "IS_RSTALLCARRYIN_INVERTED" *)
    input RSTALLCARRYIN;
    (* invertible_pin = "IS_RSTALUMODE_INVERTED" *)
    input RSTALUMODE;
    (* invertible_pin = "IS_RSTB_INVERTED" *)
    input RSTB;
    (* invertible_pin = "IS_RSTC_INVERTED" *)
    input RSTC;
    (* invertible_pin = "IS_RSTCTRL_INVERTED" *)
    input RSTCTRL;
    (* invertible_pin = "IS_RSTD_INVERTED" *)
    input RSTD;
    (* invertible_pin = "IS_RSTINMODE_INVERTED" *)
    input RSTINMODE;
    (* invertible_pin = "IS_RSTM_INVERTED" *)
    input RSTM;
    (* invertible_pin = "IS_RSTP_INVERTED" *)
    input RSTP;
endmodule

module IDELAYE2 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "IDATAIN";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter IDELAY_TYPE = "FIXED";
    parameter integer IDELAY_VALUE = 0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_DATAIN_INVERTED = 1'b0;
    parameter [0:0] IS_IDATAIN_INVERTED = 1'b0;
    parameter PIPE_SEL = "FALSE";
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    parameter integer SIM_DELAY_D = 0;
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    input CINVCTRL;
    input [4:0] CNTVALUEIN;
    (* invertible_pin = "IS_DATAIN_INVERTED" *)
    input DATAIN;
    (* invertible_pin = "IS_IDATAIN_INVERTED" *)
    input IDATAIN;
    input INC;
    input LD;
    input LDPIPEEN;
    input REGRST;
endmodule

module ODELAYE2 (...);
    parameter CINVCTRL_SEL = "FALSE";
    parameter DELAY_SRC = "ODATAIN";
    parameter HIGH_PERFORMANCE_MODE = "FALSE";
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_ODATAIN_INVERTED = 1'b0;
    parameter ODELAY_TYPE = "FIXED";
    parameter integer ODELAY_VALUE = 0;
    parameter PIPE_SEL = "FALSE";
    parameter real REFCLK_FREQUENCY = 200.0;
    parameter SIGNAL_PATTERN = "DATA";
    parameter integer SIM_DELAY_D = 0;
    output [4:0] CNTVALUEOUT;
    output DATAOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    input CE;
    input CINVCTRL;
    input CLKIN;
    input [4:0] CNTVALUEIN;
    input INC;
    input LD;
    input LDPIPEEN;
    (* invertible_pin = "IS_ODATAIN_INVERTED" *)
    input ODATAIN;
    input REGRST;
endmodule

module ISERDESE2 (...);
    parameter DATA_RATE = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter DYN_CLKDIV_INV_EN = "FALSE";
    parameter DYN_CLK_INV_EN = "FALSE";
    parameter [0:0] INIT_Q1 = 1'b0;
    parameter [0:0] INIT_Q2 = 1'b0;
    parameter [0:0] INIT_Q3 = 1'b0;
    parameter [0:0] INIT_Q4 = 1'b0;
    parameter INTERFACE_TYPE = "MEMORY";
    parameter IOBDELAY = "NONE";
    parameter [0:0] IS_CLKB_INVERTED = 1'b0;
    parameter [0:0] IS_CLKDIVP_INVERTED = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_D_INVERTED = 1'b0;
    parameter [0:0] IS_OCLKB_INVERTED = 1'b0;
    parameter [0:0] IS_OCLK_INVERTED = 1'b0;
    parameter integer NUM_CE = 2;
    parameter OFB_USED = "FALSE";
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_Q1 = 1'b0;
    parameter [0:0] SRVAL_Q2 = 1'b0;
    parameter [0:0] SRVAL_Q3 = 1'b0;
    parameter [0:0] SRVAL_Q4 = 1'b0;
    output O;
    output Q1;
    output Q2;
    output Q3;
    output Q4;
    output Q5;
    output Q6;
    output Q7;
    output Q8;
    output SHIFTOUT1;
    output SHIFTOUT2;
    input BITSLIP;
    input CE1;
    input CE2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKB_INVERTED" *)
    input CLKB;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIVP_INVERTED" *)
    input CLKDIVP;
    (* invertible_pin = "IS_D_INVERTED" *)
    input D;
    input DDLY;
    input DYNCLKDIVSEL;
    input DYNCLKSEL;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_OCLK_INVERTED" *)
    input OCLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_OCLKB_INVERTED" *)
    input OCLKB;
    input OFB;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
endmodule

module OSERDESE2 (...);
    parameter DATA_RATE_OQ = "DDR";
    parameter DATA_RATE_TQ = "DDR";
    parameter integer DATA_WIDTH = 4;
    parameter [0:0] INIT_OQ = 1'b0;
    parameter [0:0] INIT_TQ = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter [0:0] IS_D3_INVERTED = 1'b0;
    parameter [0:0] IS_D4_INVERTED = 1'b0;
    parameter [0:0] IS_D5_INVERTED = 1'b0;
    parameter [0:0] IS_D6_INVERTED = 1'b0;
    parameter [0:0] IS_D7_INVERTED = 1'b0;
    parameter [0:0] IS_D8_INVERTED = 1'b0;
    parameter [0:0] IS_T1_INVERTED = 1'b0;
    parameter [0:0] IS_T2_INVERTED = 1'b0;
    parameter [0:0] IS_T3_INVERTED = 1'b0;
    parameter [0:0] IS_T4_INVERTED = 1'b0;
    parameter SERDES_MODE = "MASTER";
    parameter [0:0] SRVAL_OQ = 1'b0;
    parameter [0:0] SRVAL_TQ = 1'b0;
    parameter TBYTE_CTL = "FALSE";
    parameter TBYTE_SRC = "FALSE";
    parameter integer TRISTATE_WIDTH = 4;
    output OFB;
    output OQ;
    output SHIFTOUT1;
    output SHIFTOUT2;
    output TBYTEOUT;
    output TFB;
    output TQ;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    (* invertible_pin = "IS_D1_INVERTED" *)
    input D1;
    (* invertible_pin = "IS_D2_INVERTED" *)
    input D2;
    (* invertible_pin = "IS_D3_INVERTED" *)
    input D3;
    (* invertible_pin = "IS_D4_INVERTED" *)
    input D4;
    (* invertible_pin = "IS_D5_INVERTED" *)
    input D5;
    (* invertible_pin = "IS_D6_INVERTED" *)
    input D6;
    (* invertible_pin = "IS_D7_INVERTED" *)
    input D7;
    (* invertible_pin = "IS_D8_INVERTED" *)
    input D8;
    input OCE;
    input RST;
    input SHIFTIN1;
    input SHIFTIN2;
    (* invertible_pin = "IS_T1_INVERTED" *)
    input T1;
    (* invertible_pin = "IS_T2_INVERTED" *)
    input T2;
    (* invertible_pin = "IS_T3_INVERTED" *)
    input T3;
    (* invertible_pin = "IS_T4_INVERTED" *)
    input T4;
    input TBYTEIN;
    input TCE;
endmodule

(* keep *)
module PHASER_IN (...);
    parameter integer CLKOUT_DIV = 4;
    parameter DQS_BIAS_MODE = "FALSE";
    parameter EN_ISERDES_RST = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter FREQ_REF_DIV = "NONE";
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter integer SEL_CLK_OFFSET = 5;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output FINEOVERFLOW;
    output ICLK;
    output ICLKDIV;
    output ISERDESRST;
    output RCLK;
    output [5:0] COUNTERREADVAL;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input DIVIDERST;
    input EDGEADV;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SYNCIN;
    input SYSCLK;
    input [1:0] RANKSEL;
    input [5:0] COUNTERLOADVAL;
endmodule

(* keep *)
module PHASER_IN_PHY (...);
    parameter BURST_MODE = "FALSE";
    parameter integer CLKOUT_DIV = 4;
    parameter [0:0] DQS_AUTO_RECAL = 1'b1;
    parameter DQS_BIAS_MODE = "FALSE";
    parameter [2:0] DQS_FIND_PATTERN = 3'b001;
    parameter integer FINE_DELAY = 0;
    parameter FREQ_REF_DIV = "NONE";
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter integer SEL_CLK_OFFSET = 5;
    parameter SYNC_IN_DIV_RST = "FALSE";
    parameter WR_CYCLES = "FALSE";
    output DQSFOUND;
    output DQSOUTOFRANGE;
    output FINEOVERFLOW;
    output ICLK;
    output ICLKDIV;
    output ISERDESRST;
    output PHASELOCKED;
    output RCLK;
    output WRENABLE;
    output [5:0] COUNTERREADVAL;
    input BURSTPENDINGPHY;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input RSTDQSFIND;
    input SYNCIN;
    input SYSCLK;
    input [1:0] ENCALIBPHY;
    input [1:0] RANKSELPHY;
    input [5:0] COUNTERLOADVAL;
endmodule

(* keep *)
module PHASER_OUT (...);
    parameter integer CLKOUT_DIV = 4;
    parameter COARSE_BYPASS = "FALSE";
    parameter integer COARSE_DELAY = 0;
    parameter EN_OSERDES_RST = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OCLKDELAY_INV = "FALSE";
    parameter integer OCLK_DELAY = 0;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter [2:0] PO = 3'b000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output COARSEOVERFLOW;
    output FINEOVERFLOW;
    output OCLK;
    output OCLKDELAYED;
    output OCLKDIV;
    output OSERDESRST;
    output [8:0] COUNTERREADVAL;
    input COARSEENABLE;
    input COARSEINC;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input DIVIDERST;
    input EDGEADV;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SELFINEOCLKDELAY;
    input SYNCIN;
    input SYSCLK;
    input [8:0] COUNTERLOADVAL;
endmodule

(* keep *)
module PHASER_OUT_PHY (...);
    parameter integer CLKOUT_DIV = 4;
    parameter COARSE_BYPASS = "FALSE";
    parameter integer COARSE_DELAY = 0;
    parameter DATA_CTL_N = "FALSE";
    parameter DATA_RD_CYCLES = "FALSE";
    parameter integer FINE_DELAY = 0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real MEMREFCLK_PERIOD = 0.000;
    parameter OCLKDELAY_INV = "FALSE";
    parameter integer OCLK_DELAY = 0;
    parameter OUTPUT_CLK_SRC = "PHASE_REF";
    parameter real PHASEREFCLK_PERIOD = 0.000;
    parameter [2:0] PO = 3'b000;
    parameter real REFCLK_PERIOD = 0.000;
    parameter SYNC_IN_DIV_RST = "FALSE";
    output COARSEOVERFLOW;
    output FINEOVERFLOW;
    output OCLK;
    output OCLKDELAYED;
    output OCLKDIV;
    output OSERDESRST;
    output RDENABLE;
    output [1:0] CTSBUS;
    output [1:0] DQSBUS;
    output [1:0] DTSBUS;
    output [8:0] COUNTERREADVAL;
    input BURSTPENDINGPHY;
    input COARSEENABLE;
    input COARSEINC;
    input COUNTERLOADEN;
    input COUNTERREADEN;
    input FINEENABLE;
    input FINEINC;
    input FREQREFCLK;
    input MEMREFCLK;
    input PHASEREFCLK;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input SELFINEOCLKDELAY;
    input SYNCIN;
    input SYSCLK;
    input [1:0] ENCALIBPHY;
    input [8:0] COUNTERLOADVAL;
endmodule

(* keep *)
module PHASER_REF (...);
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    output LOCKED;
    input CLKIN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

(* keep *)
module PHY_CONTROL (...);
    parameter integer AO_TOGGLE = 0;
    parameter [3:0] AO_WRLVL_EN = 4'b0000;
    parameter BURST_MODE = "FALSE";
    parameter integer CLK_RATIO = 1;
    parameter integer CMD_OFFSET = 0;
    parameter integer CO_DURATION = 0;
    parameter DATA_CTL_A_N = "FALSE";
    parameter DATA_CTL_B_N = "FALSE";
    parameter DATA_CTL_C_N = "FALSE";
    parameter DATA_CTL_D_N = "FALSE";
    parameter DISABLE_SEQ_MATCH = "TRUE";
    parameter integer DI_DURATION = 0;
    parameter integer DO_DURATION = 0;
    parameter integer EVENTS_DELAY = 63;
    parameter integer FOUR_WINDOW_CLOCKS = 63;
    parameter MULTI_REGION = "FALSE";
    parameter PHY_COUNT_ENABLE = "FALSE";
    parameter integer RD_CMD_OFFSET_0 = 0;
    parameter integer RD_CMD_OFFSET_1 = 00;
    parameter integer RD_CMD_OFFSET_2 = 0;
    parameter integer RD_CMD_OFFSET_3 = 0;
    parameter integer RD_DURATION_0 = 0;
    parameter integer RD_DURATION_1 = 0;
    parameter integer RD_DURATION_2 = 0;
    parameter integer RD_DURATION_3 = 0;
    parameter SYNC_MODE = "FALSE";
    parameter integer WR_CMD_OFFSET_0 = 0;
    parameter integer WR_CMD_OFFSET_1 = 0;
    parameter integer WR_CMD_OFFSET_2 = 0;
    parameter integer WR_CMD_OFFSET_3 = 0;
    parameter integer WR_DURATION_0 = 0;
    parameter integer WR_DURATION_1 = 0;
    parameter integer WR_DURATION_2 = 0;
    parameter integer WR_DURATION_3 = 0;
    output PHYCTLALMOSTFULL;
    output PHYCTLEMPTY;
    output PHYCTLFULL;
    output PHYCTLREADY;
    output [1:0] INRANKA;
    output [1:0] INRANKB;
    output [1:0] INRANKC;
    output [1:0] INRANKD;
    output [1:0] PCENABLECALIB;
    output [3:0] AUXOUTPUT;
    output [3:0] INBURSTPENDING;
    output [3:0] OUTBURSTPENDING;
    input MEMREFCLK;
    input PHYCLK;
    input PHYCTLMSTREMPTY;
    input PHYCTLWRENABLE;
    input PLLLOCK;
    input READCALIBENABLE;
    input REFDLLLOCK;
    input RESET;
    input SYNCIN;
    input WRITECALIBENABLE;
    input [31:0] PHYCTLWD;
endmodule

module IDDRE1 (...);
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter [0:0] IS_CB_INVERTED = 1'b0;
    parameter [0:0] IS_C_INVERTED = 1'b0;
    output Q1;
    output Q2;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CB_INVERTED" *)
    input CB;
    input D;
    input R;
endmodule

module ODDRE1 (...);
    parameter [0:0] IS_C_INVERTED = 1'b0;
    parameter [0:0] IS_D1_INVERTED = 1'b0;
    parameter [0:0] IS_D2_INVERTED = 1'b0;
    parameter [0:0] SRVAL = 1'b0;
    output Q;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_C_INVERTED" *)
    input C;
    (* invertible_pin = "IS_D1_INVERTED" *)
    input D1;
    (* invertible_pin = "IS_D2_INVERTED" *)
    input D2;
    input SR;
endmodule

module IDELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_SRC = "IDATAIN";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input DATAIN;
    input EN_VTC;
    input IDATAIN;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module ODELAYE3 (...);
    parameter CASCADE = "NONE";
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output CASC_OUT;
    output [8:0] CNTVALUEOUT;
    output DATAOUT;
    input CASC_IN;
    input CASC_RETURN;
    input CE;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    input ODATAIN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module ISERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter DDR_CLK_EDGE = "OPPOSITE_EDGE";
    parameter FIFO_ENABLE = "FALSE";
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter IDDR_MODE = "FALSE";
    parameter [0:0] IS_CLK_B_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output FIFO_EMPTY;
    output INTERNAL_DIVCLK;
    output [7:0] Q;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    input CLKDIV;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_B_INVERTED" *)
    input CLK_B;
    input D;
    (* clkbuf_sink *)
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module OSERDESE3 (...);
    parameter integer DATA_WIDTH = 8;
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLKDIV_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter ODDR_MODE = "FALSE";
    parameter OSERDES_D_BYPASS = "FALSE";
    parameter OSERDES_T_BYPASS = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output OQ;
    output T_OUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLKDIV_INVERTED" *)
    input CLKDIV;
    input [7:0] D;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input T;
endmodule

(* keep *)
module BITSLICE_CONTROL (...);
    parameter CTRL_CLK = "EXTERNAL";
    parameter DIV_MODE = "DIV2";
    parameter EN_CLK_TO_EXT_NORTH = "DISABLE";
    parameter EN_CLK_TO_EXT_SOUTH = "DISABLE";
    parameter EN_DYN_ODLY_MODE = "FALSE";
    parameter EN_OTHER_NCLK = "FALSE";
    parameter EN_OTHER_PCLK = "FALSE";
    parameter IDLY_VT_TRACK = "TRUE";
    parameter INV_RXCLK = "FALSE";
    parameter ODLY_VT_TRACK = "TRUE";
    parameter QDLY_VT_TRACK = "TRUE";
    parameter [5:0] READ_IDLE_COUNT = 6'h00;
    parameter REFCLK_SRC = "PLLCLK";
    parameter integer ROUNDING_FACTOR = 16;
    parameter RXGATE_EXTEND = "FALSE";
    parameter RX_CLK_PHASE_N = "SHIFT_0";
    parameter RX_CLK_PHASE_P = "SHIFT_0";
    parameter RX_GATING = "DISABLE";
    parameter SELF_CALIBRATE = "ENABLE";
    parameter SERIAL_MODE = "FALSE";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter SIM_SPEEDUP = "FAST";
    parameter real SIM_VERSION = 2.0;
    parameter TX_GATING = "DISABLE";
    output CLK_TO_EXT_NORTH;
    output CLK_TO_EXT_SOUTH;
    output DLY_RDY;
    output [6:0] DYN_DCI;
    output NCLK_NIBBLE_OUT;
    output PCLK_NIBBLE_OUT;
    output [15:0] RIU_RD_DATA;
    output RIU_VALID;
    output [39:0] RX_BIT_CTRL_OUT0;
    output [39:0] RX_BIT_CTRL_OUT1;
    output [39:0] RX_BIT_CTRL_OUT2;
    output [39:0] RX_BIT_CTRL_OUT3;
    output [39:0] RX_BIT_CTRL_OUT4;
    output [39:0] RX_BIT_CTRL_OUT5;
    output [39:0] RX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT0;
    output [39:0] TX_BIT_CTRL_OUT1;
    output [39:0] TX_BIT_CTRL_OUT2;
    output [39:0] TX_BIT_CTRL_OUT3;
    output [39:0] TX_BIT_CTRL_OUT4;
    output [39:0] TX_BIT_CTRL_OUT5;
    output [39:0] TX_BIT_CTRL_OUT6;
    output [39:0] TX_BIT_CTRL_OUT_TRI;
    output VTC_RDY;
    input CLK_FROM_EXT;
    input EN_VTC;
    input NCLK_NIBBLE_IN;
    input PCLK_NIBBLE_IN;
    input [3:0] PHY_RDCS0;
    input [3:0] PHY_RDCS1;
    input [3:0] PHY_RDEN;
    input [3:0] PHY_WRCS0;
    input [3:0] PHY_WRCS1;
    input PLL_CLK;
    input REFCLK;
    input [5:0] RIU_ADDR;
    input RIU_CLK;
    input RIU_NIBBLE_SEL;
    input [15:0] RIU_WR_DATA;
    input RIU_WR_EN;
    input RST;
    input [39:0] RX_BIT_CTRL_IN0;
    input [39:0] RX_BIT_CTRL_IN1;
    input [39:0] RX_BIT_CTRL_IN2;
    input [39:0] RX_BIT_CTRL_IN3;
    input [39:0] RX_BIT_CTRL_IN4;
    input [39:0] RX_BIT_CTRL_IN5;
    input [39:0] RX_BIT_CTRL_IN6;
    input [3:0] TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN0;
    input [39:0] TX_BIT_CTRL_IN1;
    input [39:0] TX_BIT_CTRL_IN2;
    input [39:0] TX_BIT_CTRL_IN3;
    input [39:0] TX_BIT_CTRL_IN4;
    input [39:0] TX_BIT_CTRL_IN5;
    input [39:0] TX_BIT_CTRL_IN6;
    input [39:0] TX_BIT_CTRL_IN_TRI;
endmodule

(* keep *)
module RIU_OR (...);
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    output [15:0] RIU_RD_DATA;
    output RIU_RD_VALID;
    input [15:0] RIU_RD_DATA_LOW;
    input [15:0] RIU_RD_DATA_UPP;
    input RIU_RD_VALID_LOW;
    input RIU_RD_VALID_UPP;
endmodule

module RX_BITSLICE (...);
    parameter CASCADE = "TRUE";
    parameter DATA_TYPE = "NONE";
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter integer DELAY_VALUE_EXT = 0;
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] IS_CLK_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_EXT_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    parameter UPDATE_MODE_EXT = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output [8:0] CNTVALUEOUT_EXT;
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    input CE;
    input CE_EXT;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    (* invertible_pin = "IS_CLK_EXT_INVERTED" *)
    input CLK_EXT;
    input [8:0] CNTVALUEIN;
    input [8:0] CNTVALUEIN_EXT;
    input DATAIN;
    input EN_VTC;
    input EN_VTC_EXT;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input INC;
    input INC_EXT;
    input LOAD;
    input LOAD_EXT;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
    (* invertible_pin = "IS_RST_DLY_EXT_INVERTED" *)
    input RST_DLY_EXT;
    input [39:0] RX_BIT_CTRL_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module RXTX_BITSLICE (...);
    parameter FIFO_SYNC_MODE = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_RX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RX_RST_INVERTED = 1'b0;
    parameter [0:0] IS_TX_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_TX_RST_INVERTED = 1'b0;
    parameter LOOPBACK = "FALSE";
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter RX_DATA_TYPE = "NONE";
    parameter integer RX_DATA_WIDTH = 8;
    parameter RX_DELAY_FORMAT = "TIME";
    parameter RX_DELAY_TYPE = "FIXED";
    parameter integer RX_DELAY_VALUE = 0;
    parameter real RX_REFCLK_FREQUENCY = 300.0;
    parameter RX_UPDATE_MODE = "ASYNC";
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter integer TX_DATA_WIDTH = 8;
    parameter TX_DELAY_FORMAT = "TIME";
    parameter TX_DELAY_TYPE = "FIXED";
    parameter integer TX_DELAY_VALUE = 0;
    parameter TX_OUTPUT_PHASE_90 = "FALSE";
    parameter real TX_REFCLK_FREQUENCY = 300.0;
    parameter TX_UPDATE_MODE = "ASYNC";
    output FIFO_EMPTY;
    output FIFO_WRCLK_OUT;
    output O;
    output [7:0] Q;
    output [39:0] RX_BIT_CTRL_OUT;
    output [8:0] RX_CNTVALUEOUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output [8:0] TX_CNTVALUEOUT;
    output T_OUT;
    input [7:0] D;
    input DATAIN;
    input FIFO_RD_CLK;
    input FIFO_RD_EN;
    input [39:0] RX_BIT_CTRL_IN;
    input RX_CE;
    (* invertible_pin = "IS_RX_CLK_INVERTED" *)
    input RX_CLK;
    input [8:0] RX_CNTVALUEIN;
    input RX_EN_VTC;
    input RX_INC;
    input RX_LOAD;
    (* invertible_pin = "IS_RX_RST_INVERTED" *)
    input RX_RST;
    (* invertible_pin = "IS_RX_RST_DLY_INVERTED" *)
    input RX_RST_DLY;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
    input TX_CE;
    (* invertible_pin = "IS_TX_CLK_INVERTED" *)
    input TX_CLK;
    input [8:0] TX_CNTVALUEIN;
    input TX_EN_VTC;
    input TX_INC;
    input TX_LOAD;
    (* invertible_pin = "IS_TX_RST_INVERTED" *)
    input TX_RST;
    (* invertible_pin = "IS_TX_RST_DLY_INVERTED" *)
    input TX_RST_DLY;
endmodule

module TX_BITSLICE (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter ENABLE_PRE_EMPHASIS = "FALSE";
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter TBYTE_CTL = "TBYTE_IN";
    parameter UPDATE_MODE = "ASYNC";
    output [8:0] CNTVALUEOUT;
    output O;
    output [39:0] RX_BIT_CTRL_OUT;
    output [39:0] TX_BIT_CTRL_OUT;
    output T_OUT;
    input CE;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input [7:0] D;
    input EN_VTC;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
    input [39:0] RX_BIT_CTRL_IN;
    input T;
    input TBYTE_IN;
    input [39:0] TX_BIT_CTRL_IN;
endmodule

module TX_BITSLICE_TRI (...);
    parameter integer DATA_WIDTH = 8;
    parameter DELAY_FORMAT = "TIME";
    parameter DELAY_TYPE = "FIXED";
    parameter integer DELAY_VALUE = 0;
    parameter [0:0] INIT = 1'b1;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter [0:0] IS_RST_DLY_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter NATIVE_ODELAY_BYPASS = "FALSE";
    parameter OUTPUT_PHASE_90 = "FALSE";
    parameter real REFCLK_FREQUENCY = 300.0;
    parameter SIM_DEVICE = "ULTRASCALE";
    parameter real SIM_VERSION = 2.0;
    parameter UPDATE_MODE = "ASYNC";
    output [39:0] BIT_CTRL_OUT;
    output [8:0] CNTVALUEOUT;
    output TRI_OUT;
    input [39:0] BIT_CTRL_IN;
    input CE;
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input [8:0] CNTVALUEIN;
    input EN_VTC;
    input INC;
    input LOAD;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    (* invertible_pin = "IS_RST_DLY_INVERTED" *)
    input RST_DLY;
endmodule

module IBUFE3 (...);
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    input IBUFDISABLE;
    input [3:0] OSC;
    input OSC_EN;
    input VREF;
endmodule

module IBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_DELAY_VALUE = "0";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IFD_DELAY_VALUE = "AUTO";
    parameter IOSTANDARD = "DEFAULT";
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module IBUFDSE3 (...);
    parameter DIFF_TERM = "FALSE";
    parameter DQS_BIAS = "FALSE";
    parameter IBUF_LOW_PWR = "TRUE";
    parameter IOSTANDARD = "DEFAULT";
    parameter USE_IBUFDISABLE = "FALSE";
    parameter integer SIM_INPUT_BUFFER_OFFSET = 0;
    output O;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
    input IBUFDISABLE;
    input [3:0] OSC;
    input [1:0] OSC_EN;
endmodule

module OBUFDS (...);
    parameter CAPACITANCE = "DONT_CARE";
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW = "SLOW";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input I;
endmodule

module OBUFDS_DPHY (...);
    parameter IOSTANDARD = "DEFAULT";
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input HSTX_I;
    input HSTX_T;
    input LPTX_I_N;
    input LPTX_I_P;
    input LPTX_T;
endmodule

module KEEPER (...);
    inout O;
endmodule

module PULLDOWN (...);
    output O;
endmodule

module PULLUP (...);
    output O;
endmodule

(* keep *)
module DCIRESET (...);
    output LOCKED;
    input RST;
endmodule

(* keep *)
module HPIO_VREF (...);
    parameter VREF_CNTR = "OFF";
    output VREF;
    input [6:0] FABRIC_VREF_TUNE;
endmodule

module BUFG (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFGCE (...);
    parameter CE_TYPE = "SYNC";
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    (* invertible_pin = "IS_I_INVERTED" *)
    input I;
endmodule

module BUFGCE_1 (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input I;
endmodule

module BUFGMUX (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_1 (...);
    parameter CLK_SEL_TYPE = "SYNC";
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_CTRL (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFGMUX_VIRTEX4 (...);
    (* clkbuf_driver *)
    output O;
    input I0;
    input I1;
    input S;
endmodule

module BUFG_GT (...);
    (* clkbuf_driver *)
    output O;
    input CE;
    input CEMASK;
    input CLR;
    input CLRMASK;
    input [2:0] DIV;
    input I;
endmodule

module BUFG_GT_SYNC (...);
    output CESYNC;
    output CLRSYNC;
    input CE;
    input CLK;
    input CLR;
endmodule

module BUFG_PS (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFGCE_DIV (...);
    parameter integer BUFGCE_DIVIDE = 1;
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    parameter [0:0] IS_CLR_INVERTED = 1'b0;
    parameter [0:0] IS_I_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    (* invertible_pin = "IS_CLR_INVERTED" *)
    input CLR;
    (* invertible_pin = "IS_I_INVERTED" *)
    input I;
endmodule

module BUFH (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIO (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFIODQS (...);
    parameter DQSMASK_ENABLE = "FALSE";
    (* clkbuf_driver *)
    output O;
    input DQSMASK;
    input I;
endmodule

module BUFR (...);
    parameter BUFR_DIVIDE = "BYPASS";
    parameter SIM_DEVICE = "7SERIES";
    (* clkbuf_driver *)
    output O;
    input CE;
    input CLR;
    input I;
endmodule

module BUFMR (...);
    (* clkbuf_driver *)
    output O;
    input I;
endmodule

module BUFMRCE (...);
    parameter CE_TYPE = "SYNC";
    parameter integer INIT_OUT = 0;
    parameter [0:0] IS_CE_INVERTED = 1'b0;
    (* clkbuf_driver *)
    output O;
    (* invertible_pin = "IS_CE_INVERTED" *)
    input CE;
    input I;
endmodule

module MMCM_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter CLOCK_HOLD = "FALSE";
    parameter COMPENSATION = "ZHOLD";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter real VCOCLK_FREQ_MAX = 1600.0;
    parameter real VCOCLK_FREQ_MIN = 600.0;
    parameter real CLKIN_FREQ_MAX = 800.0;
    parameter real CLKIN_FREQ_MIN = 10.0;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 10.0;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output DRDY;
    output LOCKED;
    output PSDONE;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    input PSCLK;
    input PSEN;
    input PSINCDEC;
    input PWRDWN;
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module MMCM_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLOCK_HOLD = "FALSE";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module MMCME2_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter COMPENSATION = "ZHOLD";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME2_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module PLLE2_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter COMPENSATION = "ZHOLD";
    parameter STARTUP_WAIT = "FALSE";
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter real VCOCLK_FREQ_MAX = 2133.000;
    parameter real VCOCLK_FREQ_MIN = 800.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 19.000;
    parameter real CLKPFD_FREQ_MAX = 550.0;
    parameter real CLKPFD_FREQ_MIN = 19.0;
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output DRDY;
    output LOCKED;
    output [15:0] DO;
    input CLKFBIN;
    input CLKIN1;
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input DCLK;
    input DEN;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
    input [15:0] DI;
    input [6:0] DADDR;
endmodule

module PLLE2_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT1;
    output CLKOUT2;
    output CLKOUT3;
    output CLKOUT4;
    output CLKOUT5;
    output LOCKED;
    input CLKFBIN;
    input CLKIN1;
    input PWRDWN;
    input RST;
endmodule

module MMCME3_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_CLKIN2_INVERTED" *)
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME3_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE3_ADV (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1335.000;
    parameter real VCOCLK_FREQ_MIN = 600.000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE3_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME4_ADV (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter CLKFBOUT_USE_FINE_PS = "FALSE";
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKIN2_PERIOD = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 10.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter CLKOUT0_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUT1_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter CLKOUT2_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT3_USE_FINE_PS = "FALSE";
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter CLKOUT4_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter CLKOUT5_USE_FINE_PS = "FALSE";
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter CLKOUT6_USE_FINE_PS = "FALSE";
    parameter real CLKPFD_FREQ_MAX = 550.000;
    parameter real CLKPFD_FREQ_MIN = 10.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN2_INVERTED = 1'b0;
    parameter [0:0] IS_CLKINSEL_INVERTED = 1'b0;
    parameter [0:0] IS_PSEN_INVERTED = 1'b0;
    parameter [0:0] IS_PSINCDEC_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter real REF_JITTER2 = 0.010;
    parameter SS_EN = "FALSE";
    parameter SS_MODE = "CENTER_HIGH";
    parameter integer SS_MOD_PERIOD = 10000;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1600.000;
    parameter real VCOCLK_FREQ_MIN = 800.000;
    parameter STARTUP_WAIT = "FALSE";
    output CDDCDONE;
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKFBSTOPPED;
    output CLKINSTOPPED;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    output PSDONE;
    input CDDCREQ;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_CLKIN2_INVERTED" *)
    input CLKIN2;
    (* invertible_pin = "IS_CLKINSEL_INVERTED" *)
    input CLKINSEL;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input PSCLK;
    (* invertible_pin = "IS_PSEN_INVERTED" *)
    input PSEN;
    (* invertible_pin = "IS_PSINCDEC_INVERTED" *)
    input PSINCDEC;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module MMCME4_BASE (...);
    parameter BANDWIDTH = "OPTIMIZED";
    parameter real CLKFBOUT_MULT_F = 5.000;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN1_PERIOD = 0.000;
    parameter real CLKOUT0_DIVIDE_F = 1.000;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter integer CLKOUT2_DIVIDE = 1;
    parameter real CLKOUT2_DUTY_CYCLE = 0.500;
    parameter real CLKOUT2_PHASE = 0.000;
    parameter integer CLKOUT3_DIVIDE = 1;
    parameter real CLKOUT3_DUTY_CYCLE = 0.500;
    parameter real CLKOUT3_PHASE = 0.000;
    parameter CLKOUT4_CASCADE = "FALSE";
    parameter integer CLKOUT4_DIVIDE = 1;
    parameter real CLKOUT4_DUTY_CYCLE = 0.500;
    parameter real CLKOUT4_PHASE = 0.000;
    parameter integer CLKOUT5_DIVIDE = 1;
    parameter real CLKOUT5_DUTY_CYCLE = 0.500;
    parameter real CLKOUT5_PHASE = 0.000;
    parameter integer CLKOUT6_DIVIDE = 1;
    parameter real CLKOUT6_DUTY_CYCLE = 0.500;
    parameter real CLKOUT6_PHASE = 0.000;
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN1_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER1 = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKFBOUTB;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUT2;
    output CLKOUT2B;
    output CLKOUT3;
    output CLKOUT3B;
    output CLKOUT4;
    output CLKOUT5;
    output CLKOUT6;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN1_INVERTED" *)
    input CLKIN1;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE4_ADV (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_FREQ_MAX = 1066.000;
    parameter real CLKIN_FREQ_MIN = 70.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter real CLKPFD_FREQ_MAX = 667.500;
    parameter real CLKPFD_FREQ_MIN = 70.000;
    parameter COMPENSATION = "AUTO";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    parameter real VCOCLK_FREQ_MAX = 1500.000;
    parameter real VCOCLK_FREQ_MIN = 750.000;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output [15:0] DO;
    output DRDY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    input [6:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module PLLE4_BASE (...);
    parameter integer CLKFBOUT_MULT = 5;
    parameter real CLKFBOUT_PHASE = 0.000;
    parameter real CLKIN_PERIOD = 0.000;
    parameter integer CLKOUT0_DIVIDE = 1;
    parameter real CLKOUT0_DUTY_CYCLE = 0.500;
    parameter real CLKOUT0_PHASE = 0.000;
    parameter integer CLKOUT1_DIVIDE = 1;
    parameter real CLKOUT1_DUTY_CYCLE = 0.500;
    parameter real CLKOUT1_PHASE = 0.000;
    parameter CLKOUTPHY_MODE = "VCO_2X";
    parameter integer DIVCLK_DIVIDE = 1;
    parameter [0:0] IS_CLKFBIN_INVERTED = 1'b0;
    parameter [0:0] IS_CLKIN_INVERTED = 1'b0;
    parameter [0:0] IS_PWRDWN_INVERTED = 1'b0;
    parameter [0:0] IS_RST_INVERTED = 1'b0;
    parameter real REF_JITTER = 0.010;
    parameter STARTUP_WAIT = "FALSE";
    output CLKFBOUT;
    output CLKOUT0;
    output CLKOUT0B;
    output CLKOUT1;
    output CLKOUT1B;
    output CLKOUTPHY;
    output LOCKED;
    (* invertible_pin = "IS_CLKFBIN_INVERTED" *)
    input CLKFBIN;
    (* invertible_pin = "IS_CLKIN_INVERTED" *)
    input CLKIN;
    input CLKOUTPHYEN;
    (* invertible_pin = "IS_PWRDWN_INVERTED" *)
    input PWRDWN;
    (* invertible_pin = "IS_RST_INVERTED" *)
    input RST;
endmodule

module IN_FIFO (...);
    parameter integer ALMOST_EMPTY_VALUE = 1;
    parameter integer ALMOST_FULL_VALUE = 1;
    parameter ARRAY_MODE = "ARRAY_MODE_4_X_8";
    parameter SYNCHRONOUS_MODE = "FALSE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output EMPTY;
    output FULL;
    output [7:0] Q0;
    output [7:0] Q1;
    output [7:0] Q2;
    output [7:0] Q3;
    output [7:0] Q4;
    output [7:0] Q5;
    output [7:0] Q6;
    output [7:0] Q7;
    output [7:0] Q8;
    output [7:0] Q9;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RESET;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [3:0] D0;
    input [3:0] D1;
    input [3:0] D2;
    input [3:0] D3;
    input [3:0] D4;
    input [3:0] D7;
    input [3:0] D8;
    input [3:0] D9;
    input [7:0] D5;
    input [7:0] D6;
endmodule

module OUT_FIFO (...);
    parameter integer ALMOST_EMPTY_VALUE = 1;
    parameter integer ALMOST_FULL_VALUE = 1;
    parameter ARRAY_MODE = "ARRAY_MODE_8_X_4";
    parameter OUTPUT_DISABLE = "FALSE";
    parameter SYNCHRONOUS_MODE = "FALSE";
    output ALMOSTEMPTY;
    output ALMOSTFULL;
    output EMPTY;
    output FULL;
    output [3:0] Q0;
    output [3:0] Q1;
    output [3:0] Q2;
    output [3:0] Q3;
    output [3:0] Q4;
    output [3:0] Q7;
    output [3:0] Q8;
    output [3:0] Q9;
    output [7:0] Q5;
    output [7:0] Q6;
    (* clkbuf_sink *)
    input RDCLK;
    input RDEN;
    input RESET;
    (* clkbuf_sink *)
    input WRCLK;
    input WREN;
    input [7:0] D0;
    input [7:0] D1;
    input [7:0] D2;
    input [7:0] D3;
    input [7:0] D4;
    input [7:0] D5;
    input [7:0] D6;
    input [7:0] D7;
    input [7:0] D8;
    input [7:0] D9;
endmodule

module HARD_SYNC (...);
    parameter [0:0] INIT = 1'b0;
    parameter [0:0] IS_CLK_INVERTED = 1'b0;
    parameter integer LATENCY = 2;
    output DOUT;
    (* clkbuf_sink *)
    (* invertible_pin = "IS_CLK_INVERTED" *)
    input CLK;
    input DIN;
endmodule

(* keep *)
module STARTUP_VIRTEX5 (...);
    output CFGCLK;
    output CFGMCLK;
    output DINSPI;
    output EOS;
    output TCKSPI;
    input CLK;
    input GSR;
    input GTS;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUP_VIRTEX6 (...);
    parameter PROG_USR = "FALSE";
    output CFGCLK;
    output CFGMCLK;
    output DINSPI;
    output EOS;
    output PREQ;
    output TCKSPI;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUPE2 (...);
    parameter PROG_USR = "FALSE";
    parameter real SIM_CCLK_FREQ = 0.0;
    output CFGCLK;
    output CFGMCLK;
    output EOS;
    output PREQ;
    input CLK;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module STARTUPE3 (...);
    parameter PROG_USR = "FALSE";
    parameter real SIM_CCLK_FREQ = 0.0;
    output CFGCLK;
    output CFGMCLK;
    output [3:0] DI;
    output EOS;
    output PREQ;
    input [3:0] DO;
    input [3:0] DTS;
    input FCSBO;
    input FCSBTS;
    input GSR;
    input GTS;
    input KEYCLEARB;
    input PACK;
    input USRCCLKO;
    input USRCCLKTS;
    input USRDONEO;
    input USRDONETS;
endmodule

(* keep *)
module CAPTURE_VIRTEX5 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTURE_VIRTEX6 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module CAPTUREE2 (...);
    parameter ONESHOT = "TRUE";
    input CAP;
    input CLK;
endmodule

(* keep *)
module ICAP_SPARTAN6 (...);
    parameter DEVICE_ID = 32'h04000093;
    parameter SIM_CFG_FILE_NAME = "NONE";
    output BUSY;
    output [15:0] O;
    input CLK;
    input CE;
    input WRITE;
    input [15:0] I;
endmodule

(* keep *)
module ICAP_VIRTEX5 (...);
    parameter ICAP_WIDTH = "X8";
    output BUSY;
    output [31:0] O;
    input CE;
    input CLK;
    input WRITE;
    input [31:0] I;
endmodule

(* keep *)
module ICAP_VIRTEX6 (...);
    parameter [31:0] DEVICE_ID = 32'h04244093;
    parameter ICAP_WIDTH = "X8";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output BUSY;
    output [31:0] O;
    input CLK;
    input CSB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module ICAPE2 (...);
    parameter [31:0] DEVICE_ID = 32'h04244093;
    parameter ICAP_WIDTH = "X32";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output [31:0] O;
    input CLK;
    input CSIB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module ICAPE3 (...);
    parameter [31:0] DEVICE_ID = 32'h03628093;
    parameter ICAP_AUTO_SWITCH = "DISABLE";
    parameter SIM_CFG_FILE_NAME = "NONE";
    output AVAIL;
    output [31:0] O;
    output PRDONE;
    output PRERROR;
    input CLK;
    input CSIB;
    input RDWRB;
    input [31:0] I;
endmodule

(* keep *)
module BSCAN_SPARTAN6 (...);
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCAN_VIRTEX5 (...);
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output SEL;
    output SHIFT;
    output TDI;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCAN_VIRTEX6 (...);
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

(* keep *)
module BSCANE2 (...);
    parameter DISABLE_JTAG = "FALSE";
    parameter integer JTAG_CHAIN = 1;
    output CAPTURE;
    output DRCK;
    output RESET;
    output RUNTEST;
    output SEL;
    output SHIFT;
    output TCK;
    output TDI;
    output TMS;
    output UPDATE;
    input TDO;
endmodule

module DNA_PORT (...);
    parameter [56:0] SIM_DNA_VALUE = 57'h0;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module DNA_PORTE2 (...);
    parameter [95:0] SIM_DNA_VALUE = 96'h000000000000000000000000;
    output DOUT;
    input CLK;
    input DIN;
    input READ;
    input SHIFT;
endmodule

module FRAME_ECC_VIRTEX6 (...);
    parameter FARSRC = "EFAR";
    parameter FRAME_RBT_IN_FILENAME = "NONE";
    output CRCERROR;
    output ECCERROR;
    output ECCERRORSINGLE;
    output SYNDROMEVALID;
    output [12:0] SYNDROME;
    output [23:0] FAR;
    output [4:0] SYNBIT;
    output [6:0] SYNWORD;
endmodule

module FRAME_ECCE2 (...);
    parameter FARSRC = "EFAR";
    parameter FRAME_RBT_IN_FILENAME = "NONE";
    output CRCERROR;
    output ECCERROR;
    output ECCERRORSINGLE;
    output SYNDROMEVALID;
    output [12:0] SYNDROME;
    output [25:0] FAR;
    output [4:0] SYNBIT;
    output [6:0] SYNWORD;
endmodule

module FRAME_ECCE3 (...);
    output CRCERROR;
    output ECCERRORNOTSINGLE;
    output ECCERRORSINGLE;
    output ENDOFFRAME;
    output ENDOFSCAN;
    output [25:0] FAR;
    input [1:0] FARSEL;
    input ICAPBOTCLK;
    input ICAPTOPCLK;
endmodule

module FRAME_ECCE4 (...);
    output CRCERROR;
    output ECCERRORNOTSINGLE;
    output ECCERRORSINGLE;
    output ENDOFFRAME;
    output ENDOFSCAN;
    output [26:0] FAR;
    input [1:0] FARSEL;
    input ICAPBOTCLK;
    input ICAPTOPCLK;
endmodule

module USR_ACCESS_VIRTEX5 (...);
    output CFGCLK;
    output [31:0] DATA;
    output DATAVALID;
endmodule

module USR_ACCESS_VIRTEX6 (...);
    output CFGCLK;
    output [31:0] DATA;
    output DATAVALID;
endmodule

module USR_ACCESSE2 (...);
    output CFGCLK;
    output DATAVALID;
    output [31:0] DATA;
endmodule

(* keep *)
module KEY_CLEAR (...);
    input KEYCLEARB;
endmodule

(* keep *)
module MASTER_JTAG (...);
    output TDO;
    input TCK;
    input TDI;
    input TMS;
endmodule

module EFUSE_USR (...);
    parameter [31:0] SIM_EFUSE_VALUE = 32'h00000000;
    output [31:0] EFUSEUSR;
endmodule

(* keep *)
module SYSMON (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0800;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter SIM_DEVICE = "VIRTEX5";
    parameter SIM_MONITOR_FILE = "design.txt";
    output BUSY;
    output DRDY;
    output EOC;
    output EOS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output OT;
    output [15:0] DO;
    output [2:0] ALM;
    output [4:0] CHANNEL;
    input CONVST;
    input CONVSTCLK;
    input DCLK;
    input DEN;
    input DWE;
    input RESET;
    input VN;
    input VP;
    input [15:0] DI;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input [6:0] DADDR;
endmodule

(* keep *)
module XADC (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0800;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter [15:0] INIT_58 = 16'h0;
    parameter [15:0] INIT_59 = 16'h0;
    parameter [15:0] INIT_5A = 16'h0;
    parameter [15:0] INIT_5B = 16'h0;
    parameter [15:0] INIT_5C = 16'h0;
    parameter [15:0] INIT_5D = 16'h0;
    parameter [15:0] INIT_5E = 16'h0;
    parameter [15:0] INIT_5F = 16'h0;
    parameter IS_CONVSTCLK_INVERTED = 1'b0;
    parameter IS_DCLK_INVERTED = 1'b0;
    parameter SIM_DEVICE = "7SERIES";
    parameter SIM_MONITOR_FILE = "design.txt";
    output BUSY;
    output DRDY;
    output EOC;
    output EOS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output OT;
    output [15:0] DO;
    output [7:0] ALM;
    output [4:0] CHANNEL;
    output [4:0] MUXADDR;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input DWE;
    input RESET;
    input VN;
    input VP;
    input [15:0] DI;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input [6:0] DADDR;
endmodule

(* keep *)
module SYSMONE1 (...);
    parameter [15:0] INIT_40 = 16'h0;
    parameter [15:0] INIT_41 = 16'h0;
    parameter [15:0] INIT_42 = 16'h0;
    parameter [15:0] INIT_43 = 16'h0;
    parameter [15:0] INIT_44 = 16'h0;
    parameter [15:0] INIT_45 = 16'h0;
    parameter [15:0] INIT_46 = 16'h0;
    parameter [15:0] INIT_47 = 16'h0;
    parameter [15:0] INIT_48 = 16'h0;
    parameter [15:0] INIT_49 = 16'h0;
    parameter [15:0] INIT_4A = 16'h0;
    parameter [15:0] INIT_4B = 16'h0;
    parameter [15:0] INIT_4C = 16'h0;
    parameter [15:0] INIT_4D = 16'h0;
    parameter [15:0] INIT_4E = 16'h0;
    parameter [15:0] INIT_4F = 16'h0;
    parameter [15:0] INIT_50 = 16'h0;
    parameter [15:0] INIT_51 = 16'h0;
    parameter [15:0] INIT_52 = 16'h0;
    parameter [15:0] INIT_53 = 16'h0;
    parameter [15:0] INIT_54 = 16'h0;
    parameter [15:0] INIT_55 = 16'h0;
    parameter [15:0] INIT_56 = 16'h0;
    parameter [15:0] INIT_57 = 16'h0;
    parameter [15:0] INIT_58 = 16'h0;
    parameter [15:0] INIT_59 = 16'h0;
    parameter [15:0] INIT_5A = 16'h0;
    parameter [15:0] INIT_5B = 16'h0;
    parameter [15:0] INIT_5C = 16'h0;
    parameter [15:0] INIT_5D = 16'h0;
    parameter [15:0] INIT_5E = 16'h0;
    parameter [15:0] INIT_5F = 16'h0;
    parameter [15:0] INIT_60 = 16'h0;
    parameter [15:0] INIT_61 = 16'h0;
    parameter [15:0] INIT_62 = 16'h0;
    parameter [15:0] INIT_63 = 16'h0;
    parameter [15:0] INIT_64 = 16'h0;
    parameter [15:0] INIT_65 = 16'h0;
    parameter [15:0] INIT_66 = 16'h0;
    parameter [15:0] INIT_67 = 16'h0;
    parameter [15:0] INIT_68 = 16'h0;
    parameter [15:0] INIT_69 = 16'h0;
    parameter [15:0] INIT_6A = 16'h0;
    parameter [15:0] INIT_6B = 16'h0;
    parameter [15:0] INIT_6C = 16'h0;
    parameter [15:0] INIT_6D = 16'h0;
    parameter [15:0] INIT_6E = 16'h0;
    parameter [15:0] INIT_6F = 16'h0;
    parameter [15:0] INIT_70 = 16'h0;
    parameter [15:0] INIT_71 = 16'h0;
    parameter [15:0] INIT_72 = 16'h0;
    parameter [15:0] INIT_73 = 16'h0;
    parameter [15:0] INIT_74 = 16'h0;
    parameter [15:0] INIT_75 = 16'h0;
    parameter [15:0] INIT_76 = 16'h0;
    parameter [15:0] INIT_77 = 16'h0;
    parameter [15:0] INIT_78 = 16'h0;
    parameter [15:0] INIT_79 = 16'h0;
    parameter [15:0] INIT_7A = 16'h0;
    parameter [15:0] INIT_7B = 16'h0;
    parameter [15:0] INIT_7C = 16'h0;
    parameter [15:0] INIT_7D = 16'h0;
    parameter [15:0] INIT_7E = 16'h0;
    parameter [15:0] INIT_7F = 16'h0;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    input [7:0] DADDR;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

(* keep *)
module SYSMONE4 (...);
    parameter [15:0] COMMON_N_SOURCE = 16'hFFFF;
    parameter [15:0] INIT_40 = 16'h0000;
    parameter [15:0] INIT_41 = 16'h0000;
    parameter [15:0] INIT_42 = 16'h0000;
    parameter [15:0] INIT_43 = 16'h0000;
    parameter [15:0] INIT_44 = 16'h0000;
    parameter [15:0] INIT_45 = 16'h0000;
    parameter [15:0] INIT_46 = 16'h0000;
    parameter [15:0] INIT_47 = 16'h0000;
    parameter [15:0] INIT_48 = 16'h0000;
    parameter [15:0] INIT_49 = 16'h0000;
    parameter [15:0] INIT_4A = 16'h0000;
    parameter [15:0] INIT_4B = 16'h0000;
    parameter [15:0] INIT_4C = 16'h0000;
    parameter [15:0] INIT_4D = 16'h0000;
    parameter [15:0] INIT_4E = 16'h0000;
    parameter [15:0] INIT_4F = 16'h0000;
    parameter [15:0] INIT_50 = 16'h0000;
    parameter [15:0] INIT_51 = 16'h0000;
    parameter [15:0] INIT_52 = 16'h0000;
    parameter [15:0] INIT_53 = 16'h0000;
    parameter [15:0] INIT_54 = 16'h0000;
    parameter [15:0] INIT_55 = 16'h0000;
    parameter [15:0] INIT_56 = 16'h0000;
    parameter [15:0] INIT_57 = 16'h0000;
    parameter [15:0] INIT_58 = 16'h0000;
    parameter [15:0] INIT_59 = 16'h0000;
    parameter [15:0] INIT_5A = 16'h0000;
    parameter [15:0] INIT_5B = 16'h0000;
    parameter [15:0] INIT_5C = 16'h0000;
    parameter [15:0] INIT_5D = 16'h0000;
    parameter [15:0] INIT_5E = 16'h0000;
    parameter [15:0] INIT_5F = 16'h0000;
    parameter [15:0] INIT_60 = 16'h0000;
    parameter [15:0] INIT_61 = 16'h0000;
    parameter [15:0] INIT_62 = 16'h0000;
    parameter [15:0] INIT_63 = 16'h0000;
    parameter [15:0] INIT_64 = 16'h0000;
    parameter [15:0] INIT_65 = 16'h0000;
    parameter [15:0] INIT_66 = 16'h0000;
    parameter [15:0] INIT_67 = 16'h0000;
    parameter [15:0] INIT_68 = 16'h0000;
    parameter [15:0] INIT_69 = 16'h0000;
    parameter [15:0] INIT_6A = 16'h0000;
    parameter [15:0] INIT_6B = 16'h0000;
    parameter [15:0] INIT_6C = 16'h0000;
    parameter [15:0] INIT_6D = 16'h0000;
    parameter [15:0] INIT_6E = 16'h0000;
    parameter [15:0] INIT_6F = 16'h0000;
    parameter [15:0] INIT_70 = 16'h0000;
    parameter [15:0] INIT_71 = 16'h0000;
    parameter [15:0] INIT_72 = 16'h0000;
    parameter [15:0] INIT_73 = 16'h0000;
    parameter [15:0] INIT_74 = 16'h0000;
    parameter [15:0] INIT_75 = 16'h0000;
    parameter [15:0] INIT_76 = 16'h0000;
    parameter [15:0] INIT_77 = 16'h0000;
    parameter [15:0] INIT_78 = 16'h0000;
    parameter [15:0] INIT_79 = 16'h0000;
    parameter [15:0] INIT_7A = 16'h0000;
    parameter [15:0] INIT_7B = 16'h0000;
    parameter [15:0] INIT_7C = 16'h0000;
    parameter [15:0] INIT_7D = 16'h0000;
    parameter [15:0] INIT_7E = 16'h0000;
    parameter [15:0] INIT_7F = 16'h0000;
    parameter [0:0] IS_CONVSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DCLK_INVERTED = 1'b0;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MONITOR_FILE = "design.txt";
    parameter integer SYSMON_VUSER0_BANK = 0;
    parameter SYSMON_VUSER0_MONITOR = "NONE";
    parameter integer SYSMON_VUSER1_BANK = 0;
    parameter SYSMON_VUSER1_MONITOR = "NONE";
    parameter integer SYSMON_VUSER2_BANK = 0;
    parameter SYSMON_VUSER2_MONITOR = "NONE";
    parameter integer SYSMON_VUSER3_BANK = 0;
    parameter SYSMON_VUSER3_MONITOR = "NONE";
    output [15:0] ADC_DATA;
    output [15:0] ALM;
    output BUSY;
    output [5:0] CHANNEL;
    output [15:0] DO;
    output DRDY;
    output EOC;
    output EOS;
    output I2C_SCLK_TS;
    output I2C_SDA_TS;
    output JTAGBUSY;
    output JTAGLOCKED;
    output JTAGMODIFIED;
    output [4:0] MUXADDR;
    output OT;
    output SMBALERT_TS;
    input CONVST;
    (* invertible_pin = "IS_CONVSTCLK_INVERTED" *)
    input CONVSTCLK;
    input [7:0] DADDR;
    (* invertible_pin = "IS_DCLK_INVERTED" *)
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input I2C_SCLK;
    input I2C_SDA;
    input RESET;
    input [15:0] VAUXN;
    input [15:0] VAUXP;
    input VN;
    input VP;
endmodule

module GTPA1_DUAL (...);
    parameter AC_CAP_DIS_0 = "TRUE";
    parameter AC_CAP_DIS_1 = "TRUE";
    parameter integer ALIGN_COMMA_WORD_0 = 1;
    parameter integer ALIGN_COMMA_WORD_1 = 1;
    parameter integer CB2_INH_CC_PERIOD_0 = 8;
    parameter integer CB2_INH_CC_PERIOD_1 = 8;
    parameter [4:0] CDR_PH_ADJ_TIME_0 = 5'b01010;
    parameter [4:0] CDR_PH_ADJ_TIME_1 = 5'b01010;
    parameter integer CHAN_BOND_1_MAX_SKEW_0 = 7;
    parameter integer CHAN_BOND_1_MAX_SKEW_1 = 7;
    parameter integer CHAN_BOND_2_MAX_SKEW_0 = 1;
    parameter integer CHAN_BOND_2_MAX_SKEW_1 = 1;
    parameter CHAN_BOND_KEEP_ALIGN_0 = "FALSE";
    parameter CHAN_BOND_KEEP_ALIGN_1 = "FALSE";
    parameter [9:0] CHAN_BOND_SEQ_1_1_0 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_2_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_0 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_3_1 = 10'b0001001010;
    parameter [9:0] CHAN_BOND_SEQ_1_4_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_1_4_1 = 10'b0110111100;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1_0 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_1_1 = 10'b0110111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_2_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_3_1 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_0 = 10'b0100111100;
    parameter [9:0] CHAN_BOND_SEQ_2_4_1 = 10'b0100111100;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE_1 = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE_0 = "FALSE";
    parameter CHAN_BOND_SEQ_2_USE_1 = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN_0 = 1;
    parameter integer CHAN_BOND_SEQ_LEN_1 = 1;
    parameter integer CLK25_DIVIDER_0 = 4;
    parameter integer CLK25_DIVIDER_1 = 4;
    parameter CLKINDC_B_0 = "TRUE";
    parameter CLKINDC_B_1 = "TRUE";
    parameter CLKRCV_TRST_0 = "TRUE";
    parameter CLKRCV_TRST_1 = "TRUE";
    parameter CLK_CORRECT_USE_0 = "TRUE";
    parameter CLK_CORRECT_USE_1 = "TRUE";
    parameter integer CLK_COR_ADJ_LEN_0 = 1;
    parameter integer CLK_COR_ADJ_LEN_1 = 1;
    parameter integer CLK_COR_DET_LEN_0 = 1;
    parameter integer CLK_COR_DET_LEN_1 = 1;
    parameter CLK_COR_INSERT_IDLE_FLAG_0 = "FALSE";
    parameter CLK_COR_INSERT_IDLE_FLAG_1 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_0 = "FALSE";
    parameter CLK_COR_KEEP_IDLE_1 = "FALSE";
    parameter integer CLK_COR_MAX_LAT_0 = 20;
    parameter integer CLK_COR_MAX_LAT_1 = 20;
    parameter integer CLK_COR_MIN_LAT_0 = 18;
    parameter integer CLK_COR_MIN_LAT_1 = 18;
    parameter CLK_COR_PRECEDENCE_0 = "TRUE";
    parameter CLK_COR_PRECEDENCE_1 = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT_0 = 0;
    parameter integer CLK_COR_REPEAT_WAIT_1 = 0;
    parameter [9:0] CLK_COR_SEQ_1_1_0 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4_1 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE_1 = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_1_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_2_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_3_1 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4_0 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_2_4_1 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_0 = 4'b1111;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE_1 = 4'b1111;
    parameter CLK_COR_SEQ_2_USE_0 = "FALSE";
    parameter CLK_COR_SEQ_2_USE_1 = "FALSE";
    parameter CLK_OUT_GTP_SEL_0 = "REFCLKPLL0";
    parameter CLK_OUT_GTP_SEL_1 = "REFCLKPLL1";
    parameter [1:0] CM_TRIM_0 = 2'b00;
    parameter [1:0] CM_TRIM_1 = 2'b00;
    parameter [9:0] COMMA_10B_ENABLE_0 = 10'b1111111111;
    parameter [9:0] COMMA_10B_ENABLE_1 = 10'b1111111111;
    parameter [3:0] COM_BURST_VAL_0 = 4'b1111;
    parameter [3:0] COM_BURST_VAL_1 = 4'b1111;
    parameter DEC_MCOMMA_DETECT_0 = "TRUE";
    parameter DEC_MCOMMA_DETECT_1 = "TRUE";
    parameter DEC_PCOMMA_DETECT_0 = "TRUE";
    parameter DEC_PCOMMA_DETECT_1 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_0 = "TRUE";
    parameter DEC_VALID_COMMA_ONLY_1 = "TRUE";
    parameter GTP_CFG_PWRUP_0 = "TRUE";
    parameter GTP_CFG_PWRUP_1 = "TRUE";
    parameter [9:0] MCOMMA_10B_VALUE_0 = 10'b1010000011;
    parameter [9:0] MCOMMA_10B_VALUE_1 = 10'b1010000011;
    parameter MCOMMA_DETECT_0 = "TRUE";
    parameter MCOMMA_DETECT_1 = "TRUE";
    parameter [2:0] OOBDETECT_THRESHOLD_0 = 3'b110;
    parameter [2:0] OOBDETECT_THRESHOLD_1 = 3'b110;
    parameter integer OOB_CLK_DIVIDER_0 = 4;
    parameter integer OOB_CLK_DIVIDER_1 = 4;
    parameter PCI_EXPRESS_MODE_0 = "FALSE";
    parameter PCI_EXPRESS_MODE_1 = "FALSE";
    parameter [9:0] PCOMMA_10B_VALUE_0 = 10'b0101111100;
    parameter [9:0] PCOMMA_10B_VALUE_1 = 10'b0101111100;
    parameter PCOMMA_DETECT_0 = "TRUE";
    parameter PCOMMA_DETECT_1 = "TRUE";
    parameter [2:0] PLLLKDET_CFG_0 = 3'b101;
    parameter [2:0] PLLLKDET_CFG_1 = 3'b101;
    parameter [23:0] PLL_COM_CFG_0 = 24'h21680A;
    parameter [23:0] PLL_COM_CFG_1 = 24'h21680A;
    parameter [7:0] PLL_CP_CFG_0 = 8'h00;
    parameter [7:0] PLL_CP_CFG_1 = 8'h00;
    parameter integer PLL_DIVSEL_FB_0 = 5;
    parameter integer PLL_DIVSEL_FB_1 = 5;
    parameter integer PLL_DIVSEL_REF_0 = 2;
    parameter integer PLL_DIVSEL_REF_1 = 2;
    parameter integer PLL_RXDIVSEL_OUT_0 = 1;
    parameter integer PLL_RXDIVSEL_OUT_1 = 1;
    parameter PLL_SATA_0 = "FALSE";
    parameter PLL_SATA_1 = "FALSE";
    parameter PLL_SOURCE_0 = "PLL0";
    parameter PLL_SOURCE_1 = "PLL0";
    parameter integer PLL_TXDIVSEL_OUT_0 = 1;
    parameter integer PLL_TXDIVSEL_OUT_1 = 1;
    parameter [26:0] PMA_CDR_SCAN_0 = 27'h6404040;
    parameter [26:0] PMA_CDR_SCAN_1 = 27'h6404040;
    parameter [35:0] PMA_COM_CFG_EAST = 36'h000008000;
    parameter [35:0] PMA_COM_CFG_WEST = 36'h00000A000;
    parameter [6:0] PMA_RXSYNC_CFG_0 = 7'h00;
    parameter [6:0] PMA_RXSYNC_CFG_1 = 7'h00;
    parameter [24:0] PMA_RX_CFG_0 = 25'h05CE048;
    parameter [24:0] PMA_RX_CFG_1 = 25'h05CE048;
    parameter [19:0] PMA_TX_CFG_0 = 20'h00082;
    parameter [19:0] PMA_TX_CFG_1 = 20'h00082;
    parameter RCV_TERM_GND_0 = "FALSE";
    parameter RCV_TERM_GND_1 = "FALSE";
    parameter RCV_TERM_VTTRX_0 = "TRUE";
    parameter RCV_TERM_VTTRX_1 = "TRUE";
    parameter [7:0] RXEQ_CFG_0 = 8'b01111011;
    parameter [7:0] RXEQ_CFG_1 = 8'b01111011;
    parameter [0:0] RXPRBSERR_LOOPBACK_0 = 1'b0;
    parameter [0:0] RXPRBSERR_LOOPBACK_1 = 1'b0;
    parameter RX_BUFFER_USE_0 = "TRUE";
    parameter RX_BUFFER_USE_1 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_0 = "TRUE";
    parameter RX_DECODE_SEQ_MATCH_1 = "TRUE";
    parameter RX_EN_IDLE_HOLD_CDR_0 = "FALSE";
    parameter RX_EN_IDLE_HOLD_CDR_1 = "FALSE";
    parameter RX_EN_IDLE_RESET_BUF_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_BUF_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_FR_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_FR_1 = "TRUE";
    parameter RX_EN_IDLE_RESET_PH_0 = "TRUE";
    parameter RX_EN_IDLE_RESET_PH_1 = "TRUE";
    parameter RX_EN_MODE_RESET_BUF_0 = "TRUE";
    parameter RX_EN_MODE_RESET_BUF_1 = "TRUE";
    parameter [3:0] RX_IDLE_HI_CNT_0 = 4'b1000;
    parameter [3:0] RX_IDLE_HI_CNT_1 = 4'b1000;
    parameter [3:0] RX_IDLE_LO_CNT_0 = 4'b0000;
    parameter [3:0] RX_IDLE_LO_CNT_1 = 4'b0000;
    parameter RX_LOSS_OF_SYNC_FSM_0 = "FALSE";
    parameter RX_LOSS_OF_SYNC_FSM_1 = "FALSE";
    parameter integer RX_LOS_INVALID_INCR_0 = 1;
    parameter integer RX_LOS_INVALID_INCR_1 = 1;
    parameter integer RX_LOS_THRESHOLD_0 = 4;
    parameter integer RX_LOS_THRESHOLD_1 = 4;
    parameter RX_SLIDE_MODE_0 = "PCS";
    parameter RX_SLIDE_MODE_1 = "PCS";
    parameter RX_STATUS_FMT_0 = "PCIE";
    parameter RX_STATUS_FMT_1 = "PCIE";
    parameter RX_XCLK_SEL_0 = "RXREC";
    parameter RX_XCLK_SEL_1 = "RXREC";
    parameter [2:0] SATA_BURST_VAL_0 = 3'b100;
    parameter [2:0] SATA_BURST_VAL_1 = 3'b100;
    parameter [2:0] SATA_IDLE_VAL_0 = 3'b011;
    parameter [2:0] SATA_IDLE_VAL_1 = 3'b011;
    parameter integer SATA_MAX_BURST_0 = 7;
    parameter integer SATA_MAX_BURST_1 = 7;
    parameter integer SATA_MAX_INIT_0 = 22;
    parameter integer SATA_MAX_INIT_1 = 22;
    parameter integer SATA_MAX_WAKE_0 = 7;
    parameter integer SATA_MAX_WAKE_1 = 7;
    parameter integer SATA_MIN_BURST_0 = 4;
    parameter integer SATA_MIN_BURST_1 = 4;
    parameter integer SATA_MIN_INIT_0 = 12;
    parameter integer SATA_MIN_INIT_1 = 12;
    parameter integer SATA_MIN_WAKE_0 = 4;
    parameter integer SATA_MIN_WAKE_1 = 4;
    parameter integer SIM_GTPRESET_SPEEDUP = 0;
    parameter SIM_RECEIVER_DETECT_PASS = "FALSE";
    parameter [2:0] SIM_REFCLK0_SOURCE = 3'b000;
    parameter [2:0] SIM_REFCLK1_SOURCE = 3'b000;
    parameter SIM_TX_ELEC_IDLE_LEVEL = "X";
    parameter SIM_VERSION = "2.0";
    parameter [4:0] TERMINATION_CTRL_0 = 5'b10100;
    parameter [4:0] TERMINATION_CTRL_1 = 5'b10100;
    parameter TERMINATION_OVRD_0 = "FALSE";
    parameter TERMINATION_OVRD_1 = "FALSE";
    parameter [11:0] TRANS_TIME_FROM_P2_0 = 12'h03C;
    parameter [11:0] TRANS_TIME_FROM_P2_1 = 12'h03C;
    parameter [7:0] TRANS_TIME_NON_P2_0 = 8'h19;
    parameter [7:0] TRANS_TIME_NON_P2_1 = 8'h19;
    parameter [9:0] TRANS_TIME_TO_P2_0 = 10'h064;
    parameter [9:0] TRANS_TIME_TO_P2_1 = 10'h064;
    parameter [31:0] TST_ATTR_0 = 32'h00000000;
    parameter [31:0] TST_ATTR_1 = 32'h00000000;
    parameter [2:0] TXRX_INVERT_0 = 3'b011;
    parameter [2:0] TXRX_INVERT_1 = 3'b011;
    parameter TX_BUFFER_USE_0 = "FALSE";
    parameter TX_BUFFER_USE_1 = "FALSE";
    parameter [13:0] TX_DETECT_RX_CFG_0 = 14'h1832;
    parameter [13:0] TX_DETECT_RX_CFG_1 = 14'h1832;
    parameter [2:0] TX_IDLE_DELAY_0 = 3'b011;
    parameter [2:0] TX_IDLE_DELAY_1 = 3'b011;
    parameter [1:0] TX_TDCC_CFG_0 = 2'b00;
    parameter [1:0] TX_TDCC_CFG_1 = 2'b00;
    parameter TX_XCLK_SEL_0 = "TXUSR";
    parameter TX_XCLK_SEL_1 = "TXUSR";
    output DRDY;
    output PHYSTATUS0;
    output PHYSTATUS1;
    output PLLLKDET0;
    output PLLLKDET1;
    output REFCLKOUT0;
    output REFCLKOUT1;
    output REFCLKPLL0;
    output REFCLKPLL1;
    output RESETDONE0;
    output RESETDONE1;
    output RXBYTEISALIGNED0;
    output RXBYTEISALIGNED1;
    output RXBYTEREALIGN0;
    output RXBYTEREALIGN1;
    output RXCHANBONDSEQ0;
    output RXCHANBONDSEQ1;
    output RXCHANISALIGNED0;
    output RXCHANISALIGNED1;
    output RXCHANREALIGN0;
    output RXCHANREALIGN1;
    output RXCOMMADET0;
    output RXCOMMADET1;
    output RXELECIDLE0;
    output RXELECIDLE1;
    output RXPRBSERR0;
    output RXPRBSERR1;
    output RXRECCLK0;
    output RXRECCLK1;
    output RXVALID0;
    output RXVALID1;
    output TXN0;
    output TXN1;
    output TXOUTCLK0;
    output TXOUTCLK1;
    output TXP0;
    output TXP1;
    output [15:0] DRPDO;
    output [1:0] GTPCLKFBEAST;
    output [1:0] GTPCLKFBWEST;
    output [1:0] GTPCLKOUT0;
    output [1:0] GTPCLKOUT1;
    output [1:0] RXLOSSOFSYNC0;
    output [1:0] RXLOSSOFSYNC1;
    output [1:0] TXBUFSTATUS0;
    output [1:0] TXBUFSTATUS1;
    output [2:0] RXBUFSTATUS0;
    output [2:0] RXBUFSTATUS1;
    output [2:0] RXCHBONDO;
    output [2:0] RXCLKCORCNT0;
    output [2:0] RXCLKCORCNT1;
    output [2:0] RXSTATUS0;
    output [2:0] RXSTATUS1;
    output [31:0] RXDATA0;
    output [31:0] RXDATA1;
    output [3:0] RXCHARISCOMMA0;
    output [3:0] RXCHARISCOMMA1;
    output [3:0] RXCHARISK0;
    output [3:0] RXCHARISK1;
    output [3:0] RXDISPERR0;
    output [3:0] RXDISPERR1;
    output [3:0] RXNOTINTABLE0;
    output [3:0] RXNOTINTABLE1;
    output [3:0] RXRUNDISP0;
    output [3:0] RXRUNDISP1;
    output [3:0] TXKERR0;
    output [3:0] TXKERR1;
    output [3:0] TXRUNDISP0;
    output [3:0] TXRUNDISP1;
    output [4:0] RCALOUTEAST;
    output [4:0] RCALOUTWEST;
    output [4:0] TSTOUT0;
    output [4:0] TSTOUT1;
    input CLK00;
    input CLK01;
    input CLK10;
    input CLK11;
    input CLKINEAST0;
    input CLKINEAST1;
    input CLKINWEST0;
    input CLKINWEST1;
    input DCLK;
    input DEN;
    input DWE;
    input GATERXELECIDLE0;
    input GATERXELECIDLE1;
    input GCLK00;
    input GCLK01;
    input GCLK10;
    input GCLK11;
    input GTPRESET0;
    input GTPRESET1;
    input IGNORESIGDET0;
    input IGNORESIGDET1;
    input INTDATAWIDTH0;
    input INTDATAWIDTH1;
    input PLLCLK00;
    input PLLCLK01;
    input PLLCLK10;
    input PLLCLK11;
    input PLLLKDETEN0;
    input PLLLKDETEN1;
    input PLLPOWERDOWN0;
    input PLLPOWERDOWN1;
    input PRBSCNTRESET0;
    input PRBSCNTRESET1;
    input REFCLKPWRDNB0;
    input REFCLKPWRDNB1;
    input RXBUFRESET0;
    input RXBUFRESET1;
    input RXCDRRESET0;
    input RXCDRRESET1;
    input RXCHBONDMASTER0;
    input RXCHBONDMASTER1;
    input RXCHBONDSLAVE0;
    input RXCHBONDSLAVE1;
    input RXCOMMADETUSE0;
    input RXCOMMADETUSE1;
    input RXDEC8B10BUSE0;
    input RXDEC8B10BUSE1;
    input RXENCHANSYNC0;
    input RXENCHANSYNC1;
    input RXENMCOMMAALIGN0;
    input RXENMCOMMAALIGN1;
    input RXENPCOMMAALIGN0;
    input RXENPCOMMAALIGN1;
    input RXENPMAPHASEALIGN0;
    input RXENPMAPHASEALIGN1;
    input RXN0;
    input RXN1;
    input RXP0;
    input RXP1;
    input RXPMASETPHASE0;
    input RXPMASETPHASE1;
    input RXPOLARITY0;
    input RXPOLARITY1;
    input RXRESET0;
    input RXRESET1;
    input RXSLIDE0;
    input RXSLIDE1;
    input RXUSRCLK0;
    input RXUSRCLK1;
    input RXUSRCLK20;
    input RXUSRCLK21;
    input TSTCLK0;
    input TSTCLK1;
    input TXCOMSTART0;
    input TXCOMSTART1;
    input TXCOMTYPE0;
    input TXCOMTYPE1;
    input TXDETECTRX0;
    input TXDETECTRX1;
    input TXELECIDLE0;
    input TXELECIDLE1;
    input TXENC8B10BUSE0;
    input TXENC8B10BUSE1;
    input TXENPMAPHASEALIGN0;
    input TXENPMAPHASEALIGN1;
    input TXINHIBIT0;
    input TXINHIBIT1;
    input TXPDOWNASYNCH0;
    input TXPDOWNASYNCH1;
    input TXPMASETPHASE0;
    input TXPMASETPHASE1;
    input TXPOLARITY0;
    input TXPOLARITY1;
    input TXPRBSFORCEERR0;
    input TXPRBSFORCEERR1;
    input TXRESET0;
    input TXRESET1;
    input TXUSRCLK0;
    input TXUSRCLK1;
    input TXUSRCLK20;
    input TXUSRCLK21;
    input USRCODEERR0;
    input USRCODEERR1;
    input [11:0] TSTIN0;
    input [11:0] TSTIN1;
    input [15:0] DI;
    input [1:0] GTPCLKFBSEL0EAST;
    input [1:0] GTPCLKFBSEL0WEST;
    input [1:0] GTPCLKFBSEL1EAST;
    input [1:0] GTPCLKFBSEL1WEST;
    input [1:0] RXDATAWIDTH0;
    input [1:0] RXDATAWIDTH1;
    input [1:0] RXEQMIX0;
    input [1:0] RXEQMIX1;
    input [1:0] RXPOWERDOWN0;
    input [1:0] RXPOWERDOWN1;
    input [1:0] TXDATAWIDTH0;
    input [1:0] TXDATAWIDTH1;
    input [1:0] TXPOWERDOWN0;
    input [1:0] TXPOWERDOWN1;
    input [2:0] LOOPBACK0;
    input [2:0] LOOPBACK1;
    input [2:0] REFSELDYPLL0;
    input [2:0] REFSELDYPLL1;
    input [2:0] RXCHBONDI;
    input [2:0] RXENPRBSTST0;
    input [2:0] RXENPRBSTST1;
    input [2:0] TXBUFDIFFCTRL0;
    input [2:0] TXBUFDIFFCTRL1;
    input [2:0] TXENPRBSTST0;
    input [2:0] TXENPRBSTST1;
    input [2:0] TXPREEMPHASIS0;
    input [2:0] TXPREEMPHASIS1;
    input [31:0] TXDATA0;
    input [31:0] TXDATA1;
    input [3:0] TXBYPASS8B10B0;
    input [3:0] TXBYPASS8B10B1;
    input [3:0] TXCHARDISPMODE0;
    input [3:0] TXCHARDISPMODE1;
    input [3:0] TXCHARDISPVAL0;
    input [3:0] TXCHARDISPVAL1;
    input [3:0] TXCHARISK0;
    input [3:0] TXCHARISK1;
    input [3:0] TXDIFFCTRL0;
    input [3:0] TXDIFFCTRL1;
    input [4:0] RCALINEAST;
    input [4:0] RCALINWEST;
    input [7:0] DADDR;
    input [7:0] GTPTEST0;
    input [7:0] GTPTEST1;
endmodule

module GTHE2_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [19:0] ADAPT_CFG0 = 20'h00C10;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [41:0] CFOK_CFG = 42'h24800040E80;
    parameter [5:0] CFOK_CFG2 = 6'b100000;
    parameter [5:0] CFOK_CFG3 = 6'b100000;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter [28:0] CPLL_CFG = 29'h00BC07DC;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 5;
    parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "TRUE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CLKRSVD0_INVERTED = 1'b0;
    parameter [0:0] IS_CLKRSVD1_INVERTED = 1'b0;
    parameter [0:0] IS_CPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DMONITORCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_SIGVALIDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] LOOPBACK_CFG = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [31:0] PMA_RSV = 32'b00000000000000000000000010000000;
    parameter [31:0] PMA_RSV2 = 32'b00011100000000000000000000001010;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [14:0] PMA_RSV4 = 15'b000000000001000;
    parameter [3:0] PMA_RSV5 = 4'b0000;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [82:0] RXCDR_CFG = 83'h0002007FE2000C208001A;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [8:0] RXDLY_LCFG = 9'h030;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00001000000000;
    parameter [17:0] RXLPM_LF_CFG = 18'b001001000000000000;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084020;
    parameter [23:0] RXPH_CFG = 24'hC00002;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] RXPI_CFG0 = 2'b00;
    parameter [1:0] RXPI_CFG1 = 2'b00;
    parameter [1:0] RXPI_CFG2 = 2'b00;
    parameter [1:0] RXPI_CFG3 = 2'b00;
    parameter [0:0] RXPI_CFG4 = 1'b0;
    parameter [0:0] RXPI_CFG5 = 1'b0;
    parameter [2:0] RXPI_CFG6 = 3'b100;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [23:0] RX_BIAS_CFG = 24'b000011000000000000010000;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_PD = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter [2:0] RX_DFE_AGC_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_AGC_CFG2 = 4'b0000;
    parameter [0:0] RX_DFE_AGC_OVRDEN = 1'b1;
    parameter [22:0] RX_DFE_GAIN_CFG = 23'h0020C0;
    parameter [11:0] RX_DFE_H2_CFG = 12'b000000000000;
    parameter [11:0] RX_DFE_H3_CFG = 12'b000001000000;
    parameter [10:0] RX_DFE_H4_CFG = 11'b00011100000;
    parameter [10:0] RX_DFE_H5_CFG = 11'b00011100000;
    parameter [10:0] RX_DFE_H6_CFG = 11'b00000100000;
    parameter [10:0] RX_DFE_H7_CFG = 11'b00000100000;
    parameter [32:0] RX_DFE_KL_CFG = 33'b000000000000000000000001100010000;
    parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_KL_LPM_KH_CFG2 = 4'b0010;
    parameter [0:0] RX_DFE_KL_LPM_KH_OVRDEN = 1'b1;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b10;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [3:0] RX_DFE_KL_LPM_KL_CFG2 = 4'b0010;
    parameter [0:0] RX_DFE_KL_LPM_KL_OVRDEN = 1'b1;
    parameter [15:0] RX_DFE_LPM_CFG = 16'h0080;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [53:0] RX_DFE_ST_CFG = 54'h00E100000C003F;
    parameter [16:0] RX_DFE_UT_CFG = 17'b00011100000000000;
    parameter [16:0] RX_DFE_VP_CFG = 17'b00011101010100011;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter integer RX_INT_DATAWIDTH = 0;
    parameter [12:0] RX_OS_CFG = 13'b0000010000000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "1.1";
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [8:0] TXDLY_LCFG = 9'h030;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter [0:0] TXOOB_CFG = 1'b0;
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084020;
    parameter [15:0] TXPH_CFG = 16'h0780;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b0;
    parameter [2:0] TXPI_CFG5 = 3'b100;
    parameter [0:0] TXPI_GREY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_PD = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter integer TX_INT_DATAWIDTH = 0;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [16:0] TX_RXDETECT_PRECHARGE_TIME = 17'h00000;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTREFCLKMONITOR;
    output PHYSTATUS;
    output RSOSINTDONE;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDFESLIDETAPSTARTED;
    output RXDFESLIDETAPSTROBEDONE;
    output RXDFESLIDETAPSTROBESTARTED;
    output RXDFESTADAPTDONE;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    output [14:0] DMONITOROUT;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] RXDATAVALID;
    output [1:0] RXHEADERVALID;
    output [1:0] RXSTARTOFSEQ;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXSTATUS;
    output [4:0] RXCHBONDO;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    output [5:0] RXHEADER;
    output [63:0] RXDATA;
    output [6:0] RXMONITOROUT;
    output [7:0] RXCHARISCOMMA;
    output [7:0] RXCHARISK;
    output [7:0] RXDISPERR;
    output [7:0] RXNOTINTABLE;
    input CFGRESET;
    (* invertible_pin = "IS_CLKRSVD0_INVERTED" *)
    input CLKRSVD0;
    (* invertible_pin = "IS_CLKRSVD1_INVERTED" *)
    input CLKRSVD1;
    (* invertible_pin = "IS_CPLLLOCKDETCLK_INVERTED" *)
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input CPLLRESET;
    input DMONFIFORESET;
    (* invertible_pin = "IS_DMONITORCLK_INVERTED" *)
    input DMONITORCLK;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input QPLLCLK;
    input QPLLREFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFECM1EN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFESLIDETAPADAPTEN;
    input RXDFESLIDETAPHOLD;
    input RXDFESLIDETAPINITOVRDEN;
    input RXDFESLIDETAPONLYADAPTEN;
    input RXDFESLIDETAPOVRDEN;
    input RXDFESLIDETAPSTROBE;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTNTRLEN;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXQPIEN;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    (* invertible_pin = "IS_SIGVALIDCLK_INVERTED" *)
    input SIGVALIDCLK;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input TXRATEMODE;
    input TXSTARTSEQ;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [13:0] RXADAPTSELTEST;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXMONITORSEL;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] CPLLREFCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [3:0] RXOSINTCFG;
    input [3:0] RXOSINTID0;
    input [3:0] TXDIFFCTRL;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input [4:0] RXCHBONDI;
    input [4:0] RXDFEAGCTRL;
    input [4:0] RXDFESLIDETAP;
    input [4:0] TXPIPPMSTEPSIZE;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [5:0] RXDFESLIDETAPID;
    input [63:0] TXDATA;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [7:0] TX8B10BBYPASS;
    input [7:0] TXCHARDISPMODE;
    input [7:0] TXCHARDISPVAL;
    input [7:0] TXCHARISK;
    input [8:0] DRPADDR;
endmodule

module GTHE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000040000001000;
    parameter [31:0] COMMON_CFG = 32'h0000001C;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_QPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] QPLL_CFG = 27'h0480181;
    parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
    parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
    parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
    parameter [9:0] QPLL_CP = 10'b0000011111;
    parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
    parameter [9:0] QPLL_FBDIV = 10'b0000000000;
    parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
    parameter [23:0] QPLL_INIT_CFG = 24'h000006;
    parameter [15:0] QPLL_LOCK_CFG = 16'h01E8;
    parameter [3:0] QPLL_LPF = 4'b1111;
    parameter integer QPLL_REFCLK_DIV = 2;
    parameter [0:0] QPLL_RP_COMP = 1'b0;
    parameter [1:0] QPLL_VTRL_RESET = 2'b00;
    parameter [1:0] RCAL_CFG = 2'b00;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "1.1";
    output DRPRDY;
    output QPLLFBCLKLOST;
    output QPLLLOCK;
    output QPLLOUTCLK;
    output QPLLOUTREFCLK;
    output QPLLREFCLKLOST;
    output REFCLKOUTMONITOR;
    output [15:0] DRPDO;
    output [15:0] PMARSVDOUT;
    output [7:0] QPLLDMONITOR;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input BGRCALOVRDENB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    (* invertible_pin = "IS_QPLLLOCKDETCLK_INVERTED" *)
    input QPLLLOCKDETCLK;
    input QPLLLOCKEN;
    input QPLLOUTRESET;
    input QPLLPD;
    input QPLLRESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] QPLLRSVD1;
    input [2:0] QPLLREFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] QPLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module GTPE2_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [19:0] ADAPT_CFG0 = 20'b00000000000000000000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [42:0] CFOK_CFG = 43'b1001001000000000000000001000000111010000000;
    parameter [6:0] CFOK_CFG2 = 7'b0100000;
    parameter [6:0] CFOK_CFG3 = 7'b0100000;
    parameter [0:0] CFOK_CFG4 = 1'b0;
    parameter [1:0] CFOK_CFG5 = 2'b00;
    parameter [3:0] CFOK_CFG6 = 4'b0000;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter [0:0] CLK_COMMON_SWING = 1'b0;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h010;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CLKRSVD0_INVERTED = 1'b0;
    parameter [0:0] IS_CLKRSVD1_INVERTED = 1'b0;
    parameter [0:0] IS_DMONITORCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_SIGVALIDCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] LOOPBACK_CFG = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [0:0] PMA_LOOPBACK_CFG = 1'b0;
    parameter [31:0] PMA_RSV = 32'h00000333;
    parameter [31:0] PMA_RSV2 = 32'h00002050;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [3:0] PMA_RSV4 = 4'b0000;
    parameter [0:0] PMA_RSV5 = 1'b0;
    parameter [0:0] PMA_RSV6 = 1'b0;
    parameter [0:0] PMA_RSV7 = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [82:0] RXCDR_CFG = 83'h0000107FE406001041010;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [8:0] RXDLY_LCFG = 9'h020;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [6:0] RXLPMRESET_TIME = 7'b0001111;
    parameter [0:0] RXLPM_BIAS_STARTUP_DISABLE = 1'b0;
    parameter [3:0] RXLPM_CFG = 4'b0110;
    parameter [0:0] RXLPM_CFG1 = 1'b0;
    parameter [0:0] RXLPM_CM_CFG = 1'b0;
    parameter [8:0] RXLPM_GC_CFG = 9'b111100010;
    parameter [2:0] RXLPM_GC_CFG2 = 3'b001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00001111110000;
    parameter [4:0] RXLPM_HF_CFG2 = 5'b01010;
    parameter [3:0] RXLPM_HF_CFG3 = 4'b0000;
    parameter [0:0] RXLPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [0:0] RXLPM_INCM_CFG = 1'b0;
    parameter [0:0] RXLPM_IPCM_CFG = 1'b0;
    parameter [17:0] RXLPM_LF_CFG = 18'b000000001111110000;
    parameter [4:0] RXLPM_LF_CFG2 = 5'b01010;
    parameter [2:0] RXLPM_OSINT_CFG = 3'b100;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter [4:0] RXOSCALRESET_TIMEOUT = 5'b00000;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084000;
    parameter [23:0] RXPH_CFG = 24'hC00002;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [2:0] RXPI_CFG0 = 3'b000;
    parameter [0:0] RXPI_CFG1 = 1'b0;
    parameter [0:0] RXPI_CFG2 = 1'b0;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [15:0] RX_BIAS_CFG = 16'b0000111100110011;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [13:0] RX_DEBUG_CFG = 14'b00000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [12:0] RX_OS_CFG = 13'b0001111110000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SATA_PLL_CFG = "VCO_3000MHZ";
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "1.0";
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [8:0] TXDLY_LCFG = 9'h020;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter [0:0] TXOOB_CFG = 1'b0;
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084000;
    parameter [15:0] TXPH_CFG = 16'h0400;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b0;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GREY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPTXN;
    output GTPTXP;
    output PHYSTATUS;
    output PMARSVDOUT0;
    output PMARSVDOUT1;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    output [14:0] DMONITOROUT;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] RXDATAVALID;
    output [1:0] RXSTARTOFSEQ;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [31:0] RXDATA;
    output [3:0] RXCHARISCOMMA;
    output [3:0] RXCHARISK;
    output [3:0] RXCHBONDO;
    output [3:0] RXDISPERR;
    output [3:0] RXNOTINTABLE;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    input CFGRESET;
    (* invertible_pin = "IS_CLKRSVD0_INVERTED" *)
    input CLKRSVD0;
    (* invertible_pin = "IS_CLKRSVD1_INVERTED" *)
    input CLKRSVD1;
    input DMONFIFORESET;
    (* invertible_pin = "IS_DMONITORCLK_INVERTED" *)
    input DMONITORCLK;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTPRXN;
    input GTPRXP;
    input GTRESETSEL;
    input GTRXRESET;
    input GTTXRESET;
    input PLL0CLK;
    input PLL0REFCLK;
    input PLL1CLK;
    input PLL1REFCLK;
    input PMARSVDIN0;
    input PMARSVDIN1;
    input PMARSVDIN2;
    input PMARSVDIN3;
    input PMARSVDIN4;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFOVRDEN;
    input RXLPMOSINTNTRLEN;
    input RXLPMRESET;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTNTRLEN;
    input RXOSINTOVRDEN;
    input RXOSINTPD;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    (* invertible_pin = "IS_SIGVALIDCLK_INVERTED" *)
    input SIGVALIDCLK;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXRATEMODE;
    input TXSTARTSEQ;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [13:0] RXADAPTSELTEST;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [31:0] TXDATA;
    input [3:0] RXCHBONDI;
    input [3:0] RXOSINTCFG;
    input [3:0] RXOSINTID0;
    input [3:0] TX8B10BBYPASS;
    input [3:0] TXCHARDISPMODE;
    input [3:0] TXCHARDISPVAL;
    input [3:0] TXCHARISK;
    input [3:0] TXDIFFCTRL;
    input [4:0] TXPIPPMSTEPSIZE;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [8:0] DRPADDR;
endmodule

module GTPE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000000000000000;
    parameter [31:0] COMMON_CFG = 32'h00000000;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK0_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK1_INVERTED = 1'b0;
    parameter [0:0] IS_PLL0LOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_PLL1LOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] PLL0_CFG = 27'h01F03DC;
    parameter [0:0] PLL0_DMON_CFG = 1'b0;
    parameter integer PLL0_FBDIV = 4;
    parameter integer PLL0_FBDIV_45 = 5;
    parameter [23:0] PLL0_INIT_CFG = 24'h00001E;
    parameter [8:0] PLL0_LOCK_CFG = 9'h1E8;
    parameter integer PLL0_REFCLK_DIV = 1;
    parameter [26:0] PLL1_CFG = 27'h01F03DC;
    parameter [0:0] PLL1_DMON_CFG = 1'b0;
    parameter integer PLL1_FBDIV = 4;
    parameter integer PLL1_FBDIV_45 = 5;
    parameter [23:0] PLL1_INIT_CFG = 24'h00001E;
    parameter [8:0] PLL1_LOCK_CFG = 9'h1E8;
    parameter integer PLL1_REFCLK_DIV = 1;
    parameter [7:0] PLL_CLKOUT_CFG = 8'b00000000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [2:0] SIM_PLL0REFCLK_SEL = 3'b001;
    parameter [2:0] SIM_PLL1REFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "1.0";
    output DRPRDY;
    output PLL0FBCLKLOST;
    output PLL0LOCK;
    output PLL0OUTCLK;
    output PLL0OUTREFCLK;
    output PLL0REFCLKLOST;
    output PLL1FBCLKLOST;
    output PLL1LOCK;
    output PLL1OUTCLK;
    output PLL1OUTREFCLK;
    output PLL1REFCLKLOST;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [15:0] DRPDO;
    output [15:0] PMARSVDOUT;
    output [7:0] DMONITOROUT;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input BGRCALOVRDENB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input GTEASTREFCLK0;
    input GTEASTREFCLK1;
    (* invertible_pin = "IS_GTGREFCLK0_INVERTED" *)
    input GTGREFCLK0;
    (* invertible_pin = "IS_GTGREFCLK1_INVERTED" *)
    input GTGREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTWESTREFCLK0;
    input GTWESTREFCLK1;
    (* invertible_pin = "IS_PLL0LOCKDETCLK_INVERTED" *)
    input PLL0LOCKDETCLK;
    input PLL0LOCKEN;
    input PLL0PD;
    input PLL0RESET;
    (* invertible_pin = "IS_PLL1LOCKDETCLK_INVERTED" *)
    input PLL1LOCKDETCLK;
    input PLL1LOCKEN;
    input PLL1PD;
    input PLL1RESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] PLLRSVD1;
    input [2:0] PLL0REFCLKSEL;
    input [2:0] PLL1REFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] PLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module GTXE2_CHANNEL (...);
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 1;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 1;
    parameter [23:0] CPLL_CFG = 24'hB007D8;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 5;
    parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [23:0] DMONITOR_CFG = 24'h000A00;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
    parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
    parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
    parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [2:0] GEARBOX_MODE = 3'b000;
    parameter [0:0] IS_CPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_RXUSRCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXPHDLYTSTCLK_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK2_INVERTED = 1'b0;
    parameter [0:0] IS_TXUSRCLK_INVERTED = 1'b0;
    parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [31:0] PMA_RSV = 32'h00000000;
    parameter [15:0] PMA_RSV2 = 16'h2050;
    parameter [1:0] PMA_RSV3 = 2'b00;
    parameter [31:0] PMA_RSV4 = 32'h00000000;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 61;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [71:0] RXCDR_CFG = 72'h0B000023FF20400020;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [5:0] RXCDR_LOCK_CFG = 6'b010101;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [8:0] RXDLY_LCFG = 9'h030;
    parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [13:0] RXLPM_HF_CFG = 14'b00000011110000;
    parameter [13:0] RXLPM_LF_CFG = 14'b00000011110000;
    parameter [6:0] RXOOB_CFG = 7'b0000110;
    parameter integer RXOUT_DIV = 2;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [23:0] RXPHDLY_CFG = 24'h084020;
    parameter [23:0] RXPH_CFG = 24'h000000;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [4:0] RXPMARESET_TIME = 5'b00011;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [11:0] RX_BIAS_CFG = 12'b000000000000;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter integer RX_CLK25_DIV = 7;
    parameter [0:0] RX_CLKMUX_PD = 1'b1;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [2:0] RX_CM_TRIM = 3'b100;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter [11:0] RX_DEBUG_CFG = 12'b000000000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [22:0] RX_DFE_GAIN_CFG = 23'h180E0F;
    parameter [11:0] RX_DFE_H2_CFG = 12'b000111100000;
    parameter [11:0] RX_DFE_H3_CFG = 12'b000111100000;
    parameter [10:0] RX_DFE_H4_CFG = 11'b00011110000;
    parameter [10:0] RX_DFE_H5_CFG = 11'b00011110000;
    parameter [12:0] RX_DFE_KL_CFG = 13'b0001111110000;
    parameter [31:0] RX_DFE_KL_CFG2 = 32'h3008E56A;
    parameter [15:0] RX_DFE_LPM_CFG = 16'h0904;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter [16:0] RX_DFE_UT_CFG = 17'b00111111000000000;
    parameter [16:0] RX_DFE_VP_CFG = 17'b00011111100000000;
    parameter [12:0] RX_DFE_XYD_CFG = 13'b0000000010000;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter integer RX_INT_DATAWIDTH = 0;
    parameter [12:0] RX_OS_CFG = 13'b0001111110000;
    parameter integer RX_SIG_VALID_DLY = 10;
    parameter RX_XCLK_SEL = "RXREC";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
    parameter SIM_VERSION = "4.0";
    parameter [4:0] TERM_RCAL_CFG = 5'b10000;
    parameter [0:0] TERM_RCAL_OVRD = 1'b0;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [31:0] TST_RSV = 32'h00000000;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [8:0] TXDLY_LCFG = 9'h030;
    parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 2;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [23:0] TXPHDLY_CFG = 24'h084020;
    parameter [15:0] TXPH_CFG = 16'h0780;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter integer TX_CLK25_DIV = 7;
    parameter [0:0] TX_CLKMUX_PD = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [4:0] TX_DEEMPH0 = 5'b00000;
    parameter [4:0] TX_DEEMPH1 = 5'b00000;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter integer TX_INT_DATAWIDTH = 0;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter TX_XCLK_SEL = "TXUSR";
    parameter [0:0] UCODEER_CLR = 1'b0;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTREFCLKMONITOR;
    output GTXTXN;
    output GTXTXP;
    output PHYSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output RXHEADERVALID;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPRBSERR;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRESETDONE;
    output RXSTARTOFSEQ;
    output RXVALID;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXGEARBOXREADY;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output [15:0] DRPDO;
    output [15:0] PCSRSVDOUT;
    output [1:0] RXCLKCORCNT;
    output [1:0] TXBUFSTATUS;
    output [2:0] RXBUFSTATUS;
    output [2:0] RXHEADER;
    output [2:0] RXSTATUS;
    output [4:0] RXCHBONDO;
    output [4:0] RXPHMONITOR;
    output [4:0] RXPHSLIPMONITOR;
    output [63:0] RXDATA;
    output [6:0] RXMONITOROUT;
    output [7:0] DMONITOROUT;
    output [7:0] RXCHARISCOMMA;
    output [7:0] RXCHARISK;
    output [7:0] RXDISPERR;
    output [7:0] RXNOTINTABLE;
    output [9:0] TSTOUT;
    input CFGRESET;
    (* invertible_pin = "IS_CPLLLOCKDETCLK_INVERTED" *)
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input CPLLRESET;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTXRXN;
    input GTXRXP;
    input QPLLCLK;
    input QPLLREFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input RXDDIEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFECM1EN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDFEXYDHOLD;
    input RXDFEXYDOVRDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input RXGEARBOXSLIP;
    input RXLPMEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXMCOMMAALIGNEN;
    input RXOOBRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input RXQPIEN;
    input RXSLIDE;
    input RXUSERRDY;
    (* invertible_pin = "IS_RXUSRCLK2_INVERTED" *)
    input RXUSRCLK2;
    (* invertible_pin = "IS_RXUSRCLK_INVERTED" *)
    input RXUSRCLK;
    input SETERRSTATUS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input TXDEEMPH;
    input TXDETECTRX;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXINHIBIT;
    input TXPCSRESET;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    (* invertible_pin = "IS_TXPHDLYTSTCLK_INVERTED" *)
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPISOPD;
    input TXPMARESET;
    input TXPOLARITY;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input TXPRECURSORINV;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input TXSTARTSEQ;
    input TXSWING;
    input TXUSERRDY;
    (* invertible_pin = "IS_TXUSRCLK2_INVERTED" *)
    input TXUSRCLK2;
    (* invertible_pin = "IS_TXUSRCLK_INVERTED" *)
    input TXUSRCLK;
    input [15:0] DRPDI;
    input [15:0] GTRSVD;
    input [15:0] PCSRSVDIN;
    input [19:0] TSTIN;
    input [1:0] RXELECIDLEMODE;
    input [1:0] RXMONITORSEL;
    input [1:0] RXPD;
    input [1:0] RXSYSCLKSEL;
    input [1:0] TXPD;
    input [1:0] TXSYSCLKSEL;
    input [2:0] CPLLREFCLKSEL;
    input [2:0] LOOPBACK;
    input [2:0] RXCHBONDLEVEL;
    input [2:0] RXOUTCLKSEL;
    input [2:0] RXPRBSSEL;
    input [2:0] RXRATE;
    input [2:0] TXBUFDIFFCTRL;
    input [2:0] TXHEADER;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input [2:0] TXPRBSSEL;
    input [2:0] TXRATE;
    input [3:0] CLKRSVD;
    input [3:0] TXDIFFCTRL;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN2;
    input [4:0] PMARSVDIN;
    input [4:0] RXCHBONDI;
    input [4:0] TXPOSTCURSOR;
    input [4:0] TXPRECURSOR;
    input [63:0] TXDATA;
    input [6:0] TXMAINCURSOR;
    input [6:0] TXSEQUENCE;
    input [7:0] TX8B10BBYPASS;
    input [7:0] TXCHARDISPMODE;
    input [7:0] TXCHARDISPVAL;
    input [7:0] TXCHARISK;
    input [8:0] DRPADDR;
endmodule

module GTXE2_COMMON (...);
    parameter [63:0] BIAS_CFG = 64'h0000040000001000;
    parameter [31:0] COMMON_CFG = 32'h00000000;
    parameter [0:0] IS_DRPCLK_INVERTED = 1'b0;
    parameter [0:0] IS_GTGREFCLK_INVERTED = 1'b0;
    parameter [0:0] IS_QPLLLOCKDETCLK_INVERTED = 1'b0;
    parameter [26:0] QPLL_CFG = 27'h0680181;
    parameter [3:0] QPLL_CLKOUT_CFG = 4'b0000;
    parameter [5:0] QPLL_COARSE_FREQ_OVRD = 6'b010000;
    parameter [0:0] QPLL_COARSE_FREQ_OVRD_EN = 1'b0;
    parameter [9:0] QPLL_CP = 10'b0000011111;
    parameter [0:0] QPLL_CP_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_DMONITOR_SEL = 1'b0;
    parameter [9:0] QPLL_FBDIV = 10'b0000000000;
    parameter [0:0] QPLL_FBDIV_MONITOR_EN = 1'b0;
    parameter [0:0] QPLL_FBDIV_RATIO = 1'b0;
    parameter [23:0] QPLL_INIT_CFG = 24'h000006;
    parameter [15:0] QPLL_LOCK_CFG = 16'h21E8;
    parameter [3:0] QPLL_LPF = 4'b1111;
    parameter integer QPLL_REFCLK_DIV = 2;
    parameter [2:0] SIM_QPLLREFCLK_SEL = 3'b001;
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_VERSION = "4.0";
    output DRPRDY;
    output QPLLFBCLKLOST;
    output QPLLLOCK;
    output QPLLOUTCLK;
    output QPLLOUTREFCLK;
    output QPLLREFCLKLOST;
    output REFCLKOUTMONITOR;
    output [15:0] DRPDO;
    output [7:0] QPLLDMONITOR;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    (* invertible_pin = "IS_DRPCLK_INVERTED" *)
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    (* invertible_pin = "IS_GTGREFCLK_INVERTED" *)
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    (* invertible_pin = "IS_QPLLLOCKDETCLK_INVERTED" *)
    input QPLLLOCKDETCLK;
    input QPLLLOCKEN;
    input QPLLOUTRESET;
    input QPLLPD;
    input QPLLRESET;
    input RCALENB;
    input [15:0] DRPDI;
    input [15:0] QPLLRSVD1;
    input [2:0] QPLLREFCLKSEL;
    input [4:0] BGRCALOVRD;
    input [4:0] QPLLRSVD2;
    input [7:0] DRPADDR;
    input [7:0] PMARSVD;
endmodule

module IBUFDS_GTE2 (...);
    parameter CLKCM_CFG = "TRUE";
    parameter CLKRCV_TRST = "TRUE";
    parameter CLKSWING_CFG = "TRUE";
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module GTHE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'hF800;
    parameter [15:0] ADAPT_CFG1 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0080;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h07E6;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0000;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h5080;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h07E0;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h7C42;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h4000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0060;
    parameter [15:0] RXCFOK_CFG2 = 16'h000E;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0032;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_CFG0 = 16'h0A00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h7840;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h2000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h8000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_VP_CFG0 = 16'hAA00;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0033;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "Sigcfg_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h8000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0002;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h6622;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] RXPI_CFG0 = 2'b00;
    parameter [1:0] RXPI_CFG1 = 2'b00;
    parameter [1:0] RXPI_CFG2 = 2'b00;
    parameter [1:0] RXPI_CFG3 = 2'b00;
    parameter [0:0] RXPI_CFG4 = 1'b0;
    parameter [0:0] RXPI_CFG5 = 1'b1;
    parameter [2:0] RXPI_CFG6 = 3'b000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h0AD4;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter [1:0] RX_CM_SEL = 2'b11;
    parameter [3:0] RX_CM_TRIM = 4'b0100;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [3:0] RX_DFELPM_CFG0 = 4'b0110;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter [2:0] RX_DFE_AGC_CFG1 = 3'b100;
    parameter [1:0] RX_DFE_KL_LPM_KH_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KH_CFG1 = 3'b010;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 4.0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [1:0] RX_SUM_RES_CTRL = 2'b00;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b000;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [0:0] RX_WIDEMODE_CDR = 1'b0;
    parameter RX_XCLK_SEL = "RXDES";
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATUR_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter [3:0] TXDRVBIAS_P = 4'b1100;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0980;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 4.0;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter [2:0] TX_RXDETECT_REF = 3'b100;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [1:0] WB_MODE = 2'b00;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [11:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input [2:0] LOOPBACK;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDEEMPH;
    input TXDETECTRX;
    input [3:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPOSTCURSORINV;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPRECURSORINV;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPISTRONGPDOWN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE3_COMMON (...);
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] QPLL0_CFG0 = 16'h3018;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0000;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0009;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h01E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] QPLL1_CFG0 = 16'h3018;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0000;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0000;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0009;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM0DATA1_1 = 9'b000000000;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM0_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM0_WIDTH_PIN_SEL = 1'b0;
    parameter [15:0] SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter [0:0] SDM1_DATA_PIN_SEL = 1'b0;
    parameter [0:0] SDM1_WIDTH_PIN_SEL = 1'b0;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [8:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
endmodule

module GTYE3_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'b0000000000000000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h0000;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h0000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h20F8;
    parameter [15:0] CPLL_CFG1 = 16'hA494;
    parameter [15:0] CPLL_CFG2 = 16'hF001;
    parameter [5:0] CPLL_CFG3 = 6'h00;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [7:0] CPLL_INIT_CFG1 = 8'h00;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DFE_D_X_REL_POS = 1'b0;
    parameter [0:0] DFE_VCM_COMP_EN = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h000;
    parameter [9:0] ES_PMA_CFG = 10'b0000000000;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [10:0] EVODD_PHI_CFG = 11'b00000000000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] GM_BIAS_SELECT = 1'b0;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [15:0] LOOP0_CFG = 16'h0000;
    parameter [15:0] LOOP10_CFG = 16'h0000;
    parameter [15:0] LOOP11_CFG = 16'h0000;
    parameter [15:0] LOOP12_CFG = 16'h0000;
    parameter [15:0] LOOP13_CFG = 16'h0000;
    parameter [15:0] LOOP1_CFG = 16'h0000;
    parameter [15:0] LOOP2_CFG = 16'h0000;
    parameter [15:0] LOOP3_CFG = 16'h0000;
    parameter [15:0] LOOP4_CFG = 16'h0000;
    parameter [15:0] LOOP5_CFG = 16'h0000;
    parameter [15:0] LOOP6_CFG = 16'h0000;
    parameter [15:0] LOOP7_CFG = 16'h0000;
    parameter [15:0] LOOP8_CFG = 16'h0000;
    parameter [15:0] LOOP9_CFG = 16'h0000;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [2:0] PCS_RSVD1 = 3'b000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter [1:0] PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [15:0] PMA_RSV0 = 16'h0000;
    parameter [15:0] PMA_RSV1 = 16'h0000;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0000;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG1 = 16'h0300;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0300;
    parameter [15:0] RXCDR_CFG2 = 16'h0060;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0060;
    parameter [15:0] RXCDR_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG4 = 16'h0002;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h0002;
    parameter [15:0] RXCDR_CFG5 = 16'h0000;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h0000;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0001;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [1:0] RXCFOKDONE_SRC = 2'b00;
    parameter [15:0] RXCFOK_CFG0 = 16'h3E00;
    parameter [15:0] RXCFOK_CFG1 = 16'h0042;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4C00;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h1E00;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h1900;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0200;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h001F;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h0200;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0400;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000000110;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG = 16'h0100;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [15:0] RXPI_RSV0 = 16'h0000;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h1534;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 10;
    parameter [0:0] RX_CTLE1_KHKL = 1'b0;
    parameter [0:0] RX_CTLE2_KHKL = 1'b0;
    parameter [0:0] RX_CTLE3_AGC = 1'b0;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b010;
    parameter integer RX_DFELPM_CFG0 = 6;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b0;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 2;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter [2:0] RX_DFE_KL_LPM_KL_CFG1 = 3'b010;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b0;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1000;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter integer SAS_MAX_COM = 64;
    parameter integer SAS_MIN_COM = 36;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter integer SATA_MAX_BURST = 8;
    parameter integer SATA_MAX_INIT = 21;
    parameter integer SATA_MAX_WAKE = 7;
    parameter integer SATA_MIN_BURST = 4;
    parameter integer SATA_MIN_INIT = 12;
    parameter integer SATA_MIN_WAKE = 4;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter [0:0] SIM_TX_EIDLE_DRIVE_LEVEL = 1'b0;
    parameter integer SIM_VERSION = 2;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h001F;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h2020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0001;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [15:0] TXPI_RSV0 = 16'h0000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter [0:0] TX_CLKREG_PDB = 1'b0;
    parameter [2:0] TX_CLKREG_SET = 3'b000;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [5:0] TX_DCD_CFG = 6'b000010;
    parameter [0:0] TX_DCD_EN = 1'b0;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_EML_PHI_TUNE = 1'b0;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [2:0] TX_MODE_SEL = 3'b000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h7E00;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [15:0] TX_PI_CFG0 = 16'h0000;
    parameter [15:0] TX_PI_CFG1 = 16'h0000;
    parameter [0:0] TX_PI_DIV2_MODE_B = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL0 = 1'b0;
    parameter [0:0] TX_PI_SEL_QPLL1 = 1'b0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 4;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    output [2:0] BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output [2:0] BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [16:0] DMONITOROUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [7:0] PINRSRVDAS;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output [6:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input ELPCALDVORWREN;
    input ELPCALPAORWREN;
    input EVODDPHICALDONE;
    input EVODDPHICALSTART;
    input EVODDPHIDRDEN;
    input EVODDPHIDWREN;
    input EVODDPHIXRDEN;
    input EVODDPHIXWREN;
    input EYESCANMODE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input GTRESETSEL;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTYRXN;
    input GTYRXP;
    input [2:0] LOOPBACK;
    input [15:0] LOOPRSVD;
    input LPBKRXTXSEREN;
    input LPBKTXRXSEREN;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input [4:0] PCSRSVDIN2;
    input [4:0] PMARSVDIN;
    input QPLL0CLK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RSTCLKENTX;
    input RX8B10BEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCDRRESETRSV;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input RXCOMMADETEN;
    input RXDCCFORCESTART;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEVSEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input [3:0] RXOSINTCFG;
    input RXOSINTEN;
    input RXOSINTHOLD;
    input RXOSINTOVRDEN;
    input RXOSINTSTROBE;
    input RXOSINTTESTOVRDEN;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input [2:0] TXBUFDIFFCTRL;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDIFFPD;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input TXELFORCESTART;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE3_COMMON (...);
    parameter [15:0] A_SDM1DATA1_0 = 16'b0000000000000000;
    parameter [8:0] A_SDM1DATA1_1 = 9'b000000000;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [9:0] BIAS_CFG_RSVD = 10'b0000000000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0004;
    parameter [15:0] PPF0_CFG = 16'h0FFF;
    parameter [15:0] PPF1_CFG = 16'h0FFF;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h301C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0780;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0021;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1111111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter integer QPLL0_REFCLK_DIV = 2;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h301C;
    parameter [15:0] QPLL1_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0780;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0780;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0021;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1111111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter integer QPLL1_REFCLK_DIV = 2;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_EN = 1'b1;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer SIM_VERSION = 2;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0_SEL;
    output [1:0] RXRECCLK1_SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input [1:0] SDM1WIDTH;
endmodule

module IBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module OBUFDS_GTE3 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE3_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module GTHE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter [0:0] CAPBYPASS_FORCE = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter [15:0] CKCAL_RSVD0 = 16'h4000;
    parameter [15:0] CKCAL_RSVD1 = 16'h0000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter [2:0] LPBK_BIAS_CTRL = 3'b000;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter [2:0] LPBK_IND_CTRL0 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL1 = 3'b000;
    parameter [2:0] LPBK_IND_CTRL2 = 3'b000;
    parameter [3:0] LPBK_RG_CTRL = 4'b0000;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'b0000000000000000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [2:0] PROCESS_PAR = 3'b010;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [0:0] RESET_POWERSAVE_DISABLE = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0002;
    parameter [0:0] RXDFE_PWR_SAVING = 1'b0;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [0:0] RXPI_AUTO_BW_SEL_BYPASS = 1'b0;
    parameter [15:0] RXPI_CFG0 = 16'h0002;
    parameter [15:0] RXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] RXPI_LPM = 1'b0;
    parameter [1:0] RXPI_SEL_LC = 2'b00;
    parameter [1:0] RXPI_STARTCODE = 2'b00;
    parameter [0:0] RXPI_VREFSEL = 1'b0;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 12;
    parameter [7:0] RX_CTLE3_LPF = 8'b00000000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b011;
    parameter integer RX_DFELPM_CFG0 = 0;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter [1:0] RX_DFE_AGC_CFG0 = 2'b00;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 4;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [0:0] RX_DIV2_MODE_B = 1'b0;
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter [0:0] RX_EN_HI_LR = 1'b1;
    parameter [8:0] RX_EXT_RL_CTRL = 9'b000000000;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b00;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h0000;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b1001;
    parameter [3:0] RX_SUM_RESLOAD_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b1010;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b101;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [3:0] TEMPERATURE_PAR = 4'b0010;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter [3:0] TXDRVBIAS_N = 4'b1010;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG = 16'h0000;
    parameter [1:0] TXPI_CFG0 = 2'b00;
    parameter [1:0] TXPI_CFG1 = 2'b00;
    parameter [1:0] TXPI_CFG2 = 2'b00;
    parameter [0:0] TXPI_CFG3 = 1'b0;
    parameter [0:0] TXPI_CFG4 = 1'b1;
    parameter [2:0] TXPI_CFG5 = 3'b000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_LPM = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter TXPI_PPMCLK_SEL = "TXUSRCLK2";
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [0:0] TXPI_VREFSEL = 1'b0;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter integer TX_DRVMUX_CTRL = 2;
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter [15:0] TX_PHICAL_CFG2 = 16'h0000;
    parameter integer TX_PI_BIASSET = 0;
    parameter [1:0] TX_PI_IBIAS_MID = 2'b00;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0008;
    parameter integer TX_PREDRV_CTRL = 2;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [0:0] TX_SARC_LPBK_ENB = 1'b0;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTHTXN;
    output GTHTXP;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXQPISENN;
    output RXQPISENP;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXQPISENN;
    output TXQPISENP;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTHRXN;
    input GTHRXP;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input [1:0] RXDFEAGCCTRL;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input RXPHOVRDEN;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input RXQPIEN;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input TXQPIBIASEN;
    input TXQPIWEAKPUP;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTHE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [9:0] TCONGPO;
    output TCONRSVDOUT0;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input [9:0] TCONGPI;
    input TCONPOWERUP;
    input [1:0] TCONRESET;
    input [1:0] TCONRSVDIN1;
endmodule

module GTYE4_CHANNEL (...);
    parameter [0:0] ACJTAG_DEBUG_MODE = 1'b0;
    parameter [0:0] ACJTAG_MODE = 1'b0;
    parameter [0:0] ACJTAG_RESET = 1'b0;
    parameter [15:0] ADAPT_CFG0 = 16'h9200;
    parameter [15:0] ADAPT_CFG1 = 16'h801C;
    parameter [15:0] ADAPT_CFG2 = 16'h0000;
    parameter ALIGN_COMMA_DOUBLE = "FALSE";
    parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
    parameter integer ALIGN_COMMA_WORD = 1;
    parameter ALIGN_MCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
    parameter ALIGN_PCOMMA_DET = "TRUE";
    parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
    parameter [0:0] A_RXOSCALRESET = 1'b0;
    parameter [0:0] A_RXPROGDIVRESET = 1'b0;
    parameter [0:0] A_RXTERMINATION = 1'b1;
    parameter [4:0] A_TXDIFFCTRL = 5'b01100;
    parameter [0:0] A_TXPROGDIVRESET = 1'b0;
    parameter CBCC_DATA_SOURCE_SEL = "DECODED";
    parameter [0:0] CDR_SWAP_MODE_EN = 1'b0;
    parameter [0:0] CFOK_PWRSVE_EN = 1'b1;
    parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
    parameter integer CHAN_BOND_MAX_SKEW = 7;
    parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
    parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
    parameter CHAN_BOND_SEQ_2_USE = "FALSE";
    parameter integer CHAN_BOND_SEQ_LEN = 2;
    parameter [15:0] CH_HSPMUX = 16'h2424;
    parameter [15:0] CKCAL1_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL1_CFG_1 = 16'b0101000011000000;
    parameter [15:0] CKCAL1_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL1_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_0 = 16'b1100000011000000;
    parameter [15:0] CKCAL2_CFG_1 = 16'b1000000011000000;
    parameter [15:0] CKCAL2_CFG_2 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_3 = 16'b0000000000000000;
    parameter [15:0] CKCAL2_CFG_4 = 16'b0000000000000000;
    parameter CLK_CORRECT_USE = "TRUE";
    parameter CLK_COR_KEEP_IDLE = "FALSE";
    parameter integer CLK_COR_MAX_LAT = 20;
    parameter integer CLK_COR_MIN_LAT = 18;
    parameter CLK_COR_PRECEDENCE = "TRUE";
    parameter integer CLK_COR_REPEAT_WAIT = 0;
    parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
    parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
    parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
    parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
    parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
    parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
    parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
    parameter CLK_COR_SEQ_2_USE = "FALSE";
    parameter integer CLK_COR_SEQ_LEN = 2;
    parameter [15:0] CPLL_CFG0 = 16'h01FA;
    parameter [15:0] CPLL_CFG1 = 16'h24A9;
    parameter [15:0] CPLL_CFG2 = 16'h6807;
    parameter [15:0] CPLL_CFG3 = 16'h0000;
    parameter integer CPLL_FBDIV = 4;
    parameter integer CPLL_FBDIV_45 = 4;
    parameter [15:0] CPLL_INIT_CFG0 = 16'h001E;
    parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
    parameter integer CPLL_REFCLK_DIV = 1;
    parameter [2:0] CTLE3_OCAP_EXT_CTRL = 3'b000;
    parameter [0:0] CTLE3_OCAP_EXT_EN = 1'b0;
    parameter [1:0] DDI_CTRL = 2'b00;
    parameter integer DDI_REALIGN_WAIT = 15;
    parameter DEC_MCOMMA_DETECT = "TRUE";
    parameter DEC_PCOMMA_DETECT = "TRUE";
    parameter DEC_VALID_COMMA_ONLY = "TRUE";
    parameter [0:0] DELAY_ELEC = 1'b0;
    parameter [9:0] DMONITOR_CFG0 = 10'h000;
    parameter [7:0] DMONITOR_CFG1 = 8'h00;
    parameter [0:0] ES_CLK_PHASE_SEL = 1'b0;
    parameter [5:0] ES_CONTROL = 6'b000000;
    parameter ES_ERRDET_EN = "FALSE";
    parameter ES_EYE_SCAN_EN = "FALSE";
    parameter [11:0] ES_HORZ_OFFSET = 12'h800;
    parameter [4:0] ES_PRESCALE = 5'b00000;
    parameter [15:0] ES_QUALIFIER0 = 16'h0000;
    parameter [15:0] ES_QUALIFIER1 = 16'h0000;
    parameter [15:0] ES_QUALIFIER2 = 16'h0000;
    parameter [15:0] ES_QUALIFIER3 = 16'h0000;
    parameter [15:0] ES_QUALIFIER4 = 16'h0000;
    parameter [15:0] ES_QUALIFIER5 = 16'h0000;
    parameter [15:0] ES_QUALIFIER6 = 16'h0000;
    parameter [15:0] ES_QUALIFIER7 = 16'h0000;
    parameter [15:0] ES_QUALIFIER8 = 16'h0000;
    parameter [15:0] ES_QUALIFIER9 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK0 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK1 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK2 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK3 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK4 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK5 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK6 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK7 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK8 = 16'h0000;
    parameter [15:0] ES_QUAL_MASK9 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK0 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK1 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK2 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK3 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK4 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK5 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK6 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK7 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK8 = 16'h0000;
    parameter [15:0] ES_SDATA_MASK9 = 16'h0000;
    parameter integer EYESCAN_VP_RANGE = 0;
    parameter [0:0] EYE_SCAN_SWAP_EN = 1'b0;
    parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
    parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
    parameter FTS_LANE_DESKEW_EN = "FALSE";
    parameter [4:0] GEARBOX_MODE = 5'b00000;
    parameter [0:0] ISCAN_CK_PH_SEL2 = 1'b0;
    parameter [0:0] LOCAL_MASTER = 1'b0;
    parameter integer LPBK_BIAS_CTRL = 4;
    parameter [0:0] LPBK_EN_RCAL_B = 1'b0;
    parameter [3:0] LPBK_EXT_RCAL = 4'b0000;
    parameter integer LPBK_IND_CTRL0 = 5;
    parameter integer LPBK_IND_CTRL1 = 5;
    parameter integer LPBK_IND_CTRL2 = 5;
    parameter integer LPBK_RG_CTRL = 2;
    parameter [1:0] OOBDIVCTL = 2'b00;
    parameter [0:0] OOB_PWRUP = 1'b0;
    parameter PCI3_AUTO_REALIGN = "FRST_SMPL";
    parameter [0:0] PCI3_PIPE_RX_ELECIDLE = 1'b1;
    parameter [1:0] PCI3_RX_ASYNC_EBUF_BYPASS = 2'b00;
    parameter [0:0] PCI3_RX_ELECIDLE_EI2_ENABLE = 1'b0;
    parameter [5:0] PCI3_RX_ELECIDLE_H2L_COUNT = 6'b000000;
    parameter [2:0] PCI3_RX_ELECIDLE_H2L_DISABLE = 3'b000;
    parameter [5:0] PCI3_RX_ELECIDLE_HI_COUNT = 6'b000000;
    parameter [0:0] PCI3_RX_ELECIDLE_LP4_DISABLE = 1'b0;
    parameter [0:0] PCI3_RX_FIFO_DISABLE = 1'b0;
    parameter [4:0] PCIE3_CLK_COR_EMPTY_THRSH = 5'b00000;
    parameter [5:0] PCIE3_CLK_COR_FULL_THRSH = 6'b010000;
    parameter [4:0] PCIE3_CLK_COR_MAX_LAT = 5'b01000;
    parameter [4:0] PCIE3_CLK_COR_MIN_LAT = 5'b00100;
    parameter [5:0] PCIE3_CLK_COR_THRSH_TIMER = 6'b001000;
    parameter PCIE_64B_DYN_CLKSW_DIS = "FALSE";
    parameter [15:0] PCIE_BUFG_DIV_CTRL = 16'h0000;
    parameter PCIE_GEN4_64BIT_INT_EN = "FALSE";
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN12 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN3 = 2'h0;
    parameter [1:0] PCIE_PLL_SEL_MODE_GEN4 = 2'h0;
    parameter [15:0] PCIE_RXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_RXPMA_CFG = 16'h0000;
    parameter [15:0] PCIE_TXPCS_CFG_GEN3 = 16'h0000;
    parameter [15:0] PCIE_TXPMA_CFG = 16'h0000;
    parameter PCS_PCIE_EN = "FALSE";
    parameter [15:0] PCS_RSVD0 = 16'h0000;
    parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
    parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
    parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
    parameter integer PREIQ_FREQ_BST = 0;
    parameter [0:0] RATE_SW_USE_DRP = 1'b0;
    parameter [0:0] RCLK_SIPO_DLY_ENB = 1'b0;
    parameter [0:0] RCLK_SIPO_INV_EN = 1'b0;
    parameter [2:0] RTX_BUF_CML_CTRL = 3'b010;
    parameter [1:0] RTX_BUF_TERM_CTRL = 2'b00;
    parameter [4:0] RXBUFRESET_TIME = 5'b00001;
    parameter RXBUF_ADDR_MODE = "FULL";
    parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
    parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
    parameter RXBUF_EN = "TRUE";
    parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
    parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
    parameter RXBUF_RESET_ON_EIDLE = "FALSE";
    parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
    parameter integer RXBUF_THRESH_OVFLW = 0;
    parameter RXBUF_THRESH_OVRD = "FALSE";
    parameter integer RXBUF_THRESH_UNDFLW = 4;
    parameter [4:0] RXCDRFREQRESET_TIME = 5'b10000;
    parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
    parameter [15:0] RXCDR_CFG0 = 16'h0003;
    parameter [15:0] RXCDR_CFG0_GEN3 = 16'h0003;
    parameter [15:0] RXCDR_CFG1 = 16'h0000;
    parameter [15:0] RXCDR_CFG1_GEN3 = 16'h0000;
    parameter [15:0] RXCDR_CFG2 = 16'h0164;
    parameter [9:0] RXCDR_CFG2_GEN2 = 10'h164;
    parameter [15:0] RXCDR_CFG2_GEN3 = 16'h0034;
    parameter [15:0] RXCDR_CFG2_GEN4 = 16'h0034;
    parameter [15:0] RXCDR_CFG3 = 16'h0024;
    parameter [5:0] RXCDR_CFG3_GEN2 = 6'h24;
    parameter [15:0] RXCDR_CFG3_GEN3 = 16'h0024;
    parameter [15:0] RXCDR_CFG3_GEN4 = 16'h0024;
    parameter [15:0] RXCDR_CFG4 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG4_GEN3 = 16'h5CF6;
    parameter [15:0] RXCDR_CFG5 = 16'hB46B;
    parameter [15:0] RXCDR_CFG5_GEN3 = 16'h146B;
    parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
    parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
    parameter [15:0] RXCDR_LOCK_CFG0 = 16'h0040;
    parameter [15:0] RXCDR_LOCK_CFG1 = 16'h8000;
    parameter [15:0] RXCDR_LOCK_CFG2 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG3 = 16'h0000;
    parameter [15:0] RXCDR_LOCK_CFG4 = 16'h0000;
    parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
    parameter [15:0] RXCFOK_CFG0 = 16'h0000;
    parameter [15:0] RXCFOK_CFG1 = 16'h0002;
    parameter [15:0] RXCFOK_CFG2 = 16'h002D;
    parameter [15:0] RXCKCAL1_IQ_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_I_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL1_Q_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_DX_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_D_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_S_LOOP_RST_CFG = 16'h0000;
    parameter [15:0] RXCKCAL2_X_LOOP_RST_CFG = 16'h0000;
    parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
    parameter [15:0] RXDFELPM_KL_CFG0 = 16'h0000;
    parameter [15:0] RXDFELPM_KL_CFG1 = 16'h0022;
    parameter [15:0] RXDFELPM_KL_CFG2 = 16'h0100;
    parameter [15:0] RXDFE_CFG0 = 16'h4000;
    parameter [15:0] RXDFE_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_GC_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H2_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H3_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H3_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H4_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H4_CFG1 = 16'h0003;
    parameter [15:0] RXDFE_H5_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H5_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H6_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H6_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H7_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H7_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H8_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H8_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_H9_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_H9_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HA_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HA_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HB_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HB_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HC_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HC_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HD_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HD_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HE_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HE_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_HF_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_HF_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_KH_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_KH_CFG3 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_OS_CFG1 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_UT_CFG1 = 16'h0002;
    parameter [15:0] RXDFE_UT_CFG2 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG0 = 16'h0000;
    parameter [15:0] RXDFE_VP_CFG1 = 16'h0022;
    parameter [15:0] RXDLY_CFG = 16'h0010;
    parameter [15:0] RXDLY_LCFG = 16'h0030;
    parameter RXELECIDLE_CFG = "SIGCFG_4";
    parameter integer RXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter RXGEARBOX_EN = "FALSE";
    parameter [4:0] RXISCANRESET_TIME = 5'b00001;
    parameter [15:0] RXLPM_CFG = 16'h0000;
    parameter [15:0] RXLPM_GC_CFG = 16'h1000;
    parameter [15:0] RXLPM_KH_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_KH_CFG1 = 16'h0002;
    parameter [15:0] RXLPM_OS_CFG0 = 16'h0000;
    parameter [15:0] RXLPM_OS_CFG1 = 16'h0000;
    parameter [8:0] RXOOB_CFG = 9'b000110000;
    parameter RXOOB_CLK_CFG = "PMA";
    parameter [4:0] RXOSCALRESET_TIME = 5'b00011;
    parameter integer RXOUT_DIV = 4;
    parameter [4:0] RXPCSRESET_TIME = 5'b00001;
    parameter [15:0] RXPHBEACON_CFG = 16'h0000;
    parameter [15:0] RXPHDLY_CFG = 16'h2020;
    parameter [15:0] RXPHSAMP_CFG = 16'h2100;
    parameter [15:0] RXPHSLIP_CFG = 16'h9933;
    parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] RXPI_CFG0 = 16'h0102;
    parameter [15:0] RXPI_CFG1 = 16'b0000000001010100;
    parameter RXPMACLK_SEL = "DATA";
    parameter [4:0] RXPMARESET_TIME = 5'b00001;
    parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
    parameter integer RXPRBS_LINKACQ_CNT = 15;
    parameter [0:0] RXREFCLKDIV2_SEL = 1'b0;
    parameter integer RXSLIDE_AUTO_WAIT = 7;
    parameter RXSLIDE_MODE = "OFF";
    parameter [0:0] RXSYNC_MULTILANE = 1'b0;
    parameter [0:0] RXSYNC_OVRD = 1'b0;
    parameter [0:0] RXSYNC_SKIP_DA = 1'b0;
    parameter [0:0] RX_AFE_CM_EN = 1'b0;
    parameter [15:0] RX_BIAS_CFG0 = 16'h12B0;
    parameter [5:0] RX_BUFFER_CFG = 6'b000000;
    parameter [0:0] RX_CAPFF_SARC_ENB = 1'b0;
    parameter integer RX_CLK25_DIV = 8;
    parameter [0:0] RX_CLKMUX_EN = 1'b1;
    parameter [4:0] RX_CLK_SLIP_OVRD = 5'b00000;
    parameter [3:0] RX_CM_BUF_CFG = 4'b1010;
    parameter [0:0] RX_CM_BUF_PD = 1'b0;
    parameter integer RX_CM_SEL = 3;
    parameter integer RX_CM_TRIM = 12;
    parameter [0:0] RX_CTLE_PWR_SAVING = 1'b0;
    parameter [3:0] RX_CTLE_RES_CTRL = 4'b0000;
    parameter integer RX_DATA_WIDTH = 20;
    parameter [5:0] RX_DDI_SEL = 6'b000000;
    parameter RX_DEFER_RESET_BUF_EN = "TRUE";
    parameter [2:0] RX_DEGEN_CTRL = 3'b100;
    parameter integer RX_DFELPM_CFG0 = 0;
    parameter [0:0] RX_DFELPM_CFG1 = 1'b1;
    parameter [0:0] RX_DFELPM_KLKH_AGC_STUP_EN = 1'b1;
    parameter integer RX_DFE_AGC_CFG1 = 4;
    parameter integer RX_DFE_KL_LPM_KH_CFG0 = 1;
    parameter integer RX_DFE_KL_LPM_KH_CFG1 = 4;
    parameter [1:0] RX_DFE_KL_LPM_KL_CFG0 = 2'b01;
    parameter integer RX_DFE_KL_LPM_KL_CFG1 = 4;
    parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
    parameter RX_DISPERR_SEQ_MATCH = "TRUE";
    parameter [4:0] RX_DIVRESET_TIME = 5'b00001;
    parameter [0:0] RX_EN_CTLE_RCAL_B = 1'b0;
    parameter integer RX_EN_SUM_RCAL_B = 0;
    parameter [6:0] RX_EYESCAN_VS_CODE = 7'b0000000;
    parameter [0:0] RX_EYESCAN_VS_NEG_DIR = 1'b0;
    parameter [1:0] RX_EYESCAN_VS_RANGE = 2'b10;
    parameter [0:0] RX_EYESCAN_VS_UT_SIGN = 1'b0;
    parameter [0:0] RX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] RX_I2V_FILTER_EN = 1'b1;
    parameter integer RX_INT_DATAWIDTH = 1;
    parameter [0:0] RX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] RX_PMA_RSV0 = 16'h000F;
    parameter real RX_PROGDIV_CFG = 0.0;
    parameter [15:0] RX_PROGDIV_RATE = 16'h0001;
    parameter [3:0] RX_RESLOAD_CTRL = 4'b0000;
    parameter [0:0] RX_RESLOAD_OVRD = 1'b0;
    parameter [2:0] RX_SAMPLE_PERIOD = 3'b101;
    parameter integer RX_SIG_VALID_DLY = 11;
    parameter integer RX_SUM_DEGEN_AVTT_OVERITE = 0;
    parameter [0:0] RX_SUM_DFETAPREP_EN = 1'b0;
    parameter [3:0] RX_SUM_IREF_TUNE = 4'b0000;
    parameter integer RX_SUM_PWR_SAVING = 0;
    parameter [3:0] RX_SUM_RES_CTRL = 4'b0000;
    parameter [3:0] RX_SUM_VCMTUNE = 4'b0011;
    parameter [0:0] RX_SUM_VCM_BIAS_TUNE_EN = 1'b1;
    parameter [0:0] RX_SUM_VCM_OVWR = 1'b0;
    parameter [2:0] RX_SUM_VREF_TUNE = 3'b100;
    parameter [1:0] RX_TUNE_AFE_OS = 2'b00;
    parameter [2:0] RX_VREG_CTRL = 3'b010;
    parameter [0:0] RX_VREG_PDB = 1'b1;
    parameter [1:0] RX_WIDEMODE_CDR = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN3 = 2'b01;
    parameter [1:0] RX_WIDEMODE_CDR_GEN4 = 2'b01;
    parameter RX_XCLK_SEL = "RXDES";
    parameter [0:0] RX_XMODE_SEL = 1'b0;
    parameter [0:0] SAMPLE_CLK_PHASE = 1'b0;
    parameter [0:0] SAS_12G_MODE = 1'b0;
    parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
    parameter [2:0] SATA_BURST_VAL = 3'b100;
    parameter SATA_CPLL_CFG = "VCO_3000MHZ";
    parameter [2:0] SATA_EIDLE_VAL = 3'b100;
    parameter SHOW_REALIGN_COMMA = "TRUE";
    parameter SIM_MODE = "FAST";
    parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [0:0] SRSTMODE = 1'b0;
    parameter [1:0] TAPDLY_SET_TX = 2'h0;
    parameter [14:0] TERM_RCAL_CFG = 15'b100001000010000;
    parameter [2:0] TERM_RCAL_OVRD = 3'b000;
    parameter [7:0] TRANS_TIME_RATE = 8'h0E;
    parameter [7:0] TST_RSV0 = 8'h00;
    parameter [7:0] TST_RSV1 = 8'h00;
    parameter TXBUF_EN = "TRUE";
    parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
    parameter [15:0] TXDLY_CFG = 16'h0010;
    parameter [15:0] TXDLY_LCFG = 16'h0030;
    parameter integer TXDRV_FREQBAND = 0;
    parameter [15:0] TXFE_CFG0 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG1 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG2 = 16'b0000000000000000;
    parameter [15:0] TXFE_CFG3 = 16'b0000000000000000;
    parameter TXFIFO_ADDR_CFG = "LOW";
    parameter integer TXGBOX_FIFO_INIT_RD_ADDR = 4;
    parameter TXGEARBOX_EN = "FALSE";
    parameter integer TXOUT_DIV = 4;
    parameter [4:0] TXPCSRESET_TIME = 5'b00001;
    parameter [15:0] TXPHDLY_CFG0 = 16'h6020;
    parameter [15:0] TXPHDLY_CFG1 = 16'h0002;
    parameter [15:0] TXPH_CFG = 16'h0123;
    parameter [15:0] TXPH_CFG2 = 16'h0000;
    parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
    parameter [15:0] TXPI_CFG0 = 16'b0000000100000000;
    parameter [15:0] TXPI_CFG1 = 16'b0000000000000000;
    parameter [0:0] TXPI_GRAY_SEL = 1'b0;
    parameter [0:0] TXPI_INVSTROBE_SEL = 1'b0;
    parameter [0:0] TXPI_PPM = 1'b0;
    parameter [7:0] TXPI_PPM_CFG = 8'b00000000;
    parameter [2:0] TXPI_SYNFREQ_PPM = 3'b000;
    parameter [4:0] TXPMARESET_TIME = 5'b00001;
    parameter [0:0] TXREFCLKDIV2_SEL = 1'b0;
    parameter integer TXSWBST_BST = 1;
    parameter integer TXSWBST_EN = 0;
    parameter integer TXSWBST_MAG = 6;
    parameter [0:0] TXSYNC_MULTILANE = 1'b0;
    parameter [0:0] TXSYNC_OVRD = 1'b0;
    parameter [0:0] TXSYNC_SKIP_DA = 1'b0;
    parameter integer TX_CLK25_DIV = 8;
    parameter [0:0] TX_CLKMUX_EN = 1'b1;
    parameter integer TX_DATA_WIDTH = 20;
    parameter [15:0] TX_DCC_LOOP_RST_CFG = 16'h0000;
    parameter [5:0] TX_DEEMPH0 = 6'b000000;
    parameter [5:0] TX_DEEMPH1 = 6'b000000;
    parameter [5:0] TX_DEEMPH2 = 6'b000000;
    parameter [5:0] TX_DEEMPH3 = 6'b000000;
    parameter [4:0] TX_DIVRESET_TIME = 5'b00001;
    parameter TX_DRIVE_MODE = "DIRECT";
    parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
    parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
    parameter [0:0] TX_FABINT_USRCLK_FLOP = 1'b0;
    parameter [0:0] TX_FIFO_BYP_EN = 1'b0;
    parameter [0:0] TX_IDLE_DATA_ZERO = 1'b0;
    parameter integer TX_INT_DATAWIDTH = 1;
    parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
    parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
    parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
    parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
    parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
    parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
    parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
    parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
    parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
    parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
    parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
    parameter [15:0] TX_PHICAL_CFG0 = 16'h0000;
    parameter [15:0] TX_PHICAL_CFG1 = 16'h003F;
    parameter integer TX_PI_BIASSET = 0;
    parameter [0:0] TX_PMADATA_OPT = 1'b0;
    parameter [0:0] TX_PMA_POWER_SAVE = 1'b0;
    parameter [15:0] TX_PMA_RSV0 = 16'h0000;
    parameter [15:0] TX_PMA_RSV1 = 16'h0000;
    parameter TX_PROGCLK_SEL = "POSTPI";
    parameter real TX_PROGDIV_CFG = 0.0;
    parameter [15:0] TX_PROGDIV_RATE = 16'h0001;
    parameter [13:0] TX_RXDETECT_CFG = 14'h0032;
    parameter integer TX_RXDETECT_REF = 3;
    parameter [2:0] TX_SAMPLE_PERIOD = 3'b101;
    parameter [1:0] TX_SW_MEAS = 2'b00;
    parameter [2:0] TX_VREG_CTRL = 3'b000;
    parameter [0:0] TX_VREG_PDB = 1'b0;
    parameter [1:0] TX_VREG_VREFSEL = 2'b00;
    parameter TX_XCLK_SEL = "TXOUT";
    parameter [0:0] USB_BOTH_BURST_IDLE = 1'b0;
    parameter [6:0] USB_BURSTMAX_U3WAKE = 7'b1111111;
    parameter [6:0] USB_BURSTMIN_U3WAKE = 7'b1100011;
    parameter [0:0] USB_CLK_COR_EQ_EN = 1'b0;
    parameter [0:0] USB_EXT_CNTL = 1'b1;
    parameter [9:0] USB_IDLEMAX_POLLING = 10'b1010111011;
    parameter [9:0] USB_IDLEMIN_POLLING = 10'b0100101011;
    parameter [8:0] USB_LFPSPING_BURST = 9'b000000101;
    parameter [8:0] USB_LFPSPOLLING_BURST = 9'b000110001;
    parameter [8:0] USB_LFPSPOLLING_IDLE_MS = 9'b000000100;
    parameter [8:0] USB_LFPSU1EXIT_BURST = 9'b000011101;
    parameter [8:0] USB_LFPSU2LPEXIT_BURST_MS = 9'b001100011;
    parameter [8:0] USB_LFPSU3WAKE_BURST_MS = 9'b111110011;
    parameter [3:0] USB_LFPS_TPERIOD = 4'b0011;
    parameter [0:0] USB_LFPS_TPERIOD_ACCURATE = 1'b1;
    parameter [0:0] USB_MODE = 1'b0;
    parameter [0:0] USB_PCIE_ERR_REP_DIS = 1'b0;
    parameter integer USB_PING_SATA_MAX_INIT = 21;
    parameter integer USB_PING_SATA_MIN_INIT = 12;
    parameter integer USB_POLL_SATA_MAX_BURST = 8;
    parameter integer USB_POLL_SATA_MIN_BURST = 4;
    parameter [0:0] USB_RAW_ELEC = 1'b0;
    parameter [0:0] USB_RXIDLE_P0_CTRL = 1'b1;
    parameter [0:0] USB_TXIDLE_TUNE_ENABLE = 1'b1;
    parameter integer USB_U1_SATA_MAX_WAKE = 7;
    parameter integer USB_U1_SATA_MIN_WAKE = 4;
    parameter integer USB_U2_SAS_MAX_COM = 64;
    parameter integer USB_U2_SAS_MIN_COM = 36;
    parameter [0:0] USE_PCS_CLK_PHASE_SEL = 1'b0;
    parameter [0:0] Y_ALL_MODE = 1'b0;
    output BUFGTCE;
    output [2:0] BUFGTCEMASK;
    output [8:0] BUFGTDIV;
    output BUFGTRESET;
    output [2:0] BUFGTRSTMASK;
    output CPLLFBCLKLOST;
    output CPLLLOCK;
    output CPLLREFCLKLOST;
    output [15:0] DMONITOROUT;
    output DMONITOROUTCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output EYESCANDATAERROR;
    output GTPOWERGOOD;
    output GTREFCLKMONITOR;
    output GTYTXN;
    output GTYTXP;
    output PCIERATEGEN3;
    output PCIERATEIDLE;
    output [1:0] PCIERATEQPLLPD;
    output [1:0] PCIERATEQPLLRESET;
    output PCIESYNCTXSYNCDONE;
    output PCIEUSERGEN3RDY;
    output PCIEUSERPHYSTATUSRST;
    output PCIEUSERRATESTART;
    output [15:0] PCSRSVDOUT;
    output PHYSTATUS;
    output [15:0] PINRSRVDAS;
    output POWERPRESENT;
    output RESETEXCEPTION;
    output [2:0] RXBUFSTATUS;
    output RXBYTEISALIGNED;
    output RXBYTEREALIGN;
    output RXCDRLOCK;
    output RXCDRPHDONE;
    output RXCHANBONDSEQ;
    output RXCHANISALIGNED;
    output RXCHANREALIGN;
    output [4:0] RXCHBONDO;
    output RXCKCALDONE;
    output [1:0] RXCLKCORCNT;
    output RXCOMINITDET;
    output RXCOMMADET;
    output RXCOMSASDET;
    output RXCOMWAKEDET;
    output [15:0] RXCTRL0;
    output [15:0] RXCTRL1;
    output [7:0] RXCTRL2;
    output [7:0] RXCTRL3;
    output [127:0] RXDATA;
    output [7:0] RXDATAEXTENDRSVD;
    output [1:0] RXDATAVALID;
    output RXDLYSRESETDONE;
    output RXELECIDLE;
    output [5:0] RXHEADER;
    output [1:0] RXHEADERVALID;
    output RXLFPSTRESETDET;
    output RXLFPSU2LPEXITDET;
    output RXLFPSU3WAKEDET;
    output [7:0] RXMONITOROUT;
    output RXOSINTDONE;
    output RXOSINTSTARTED;
    output RXOSINTSTROBEDONE;
    output RXOSINTSTROBESTARTED;
    output RXOUTCLK;
    output RXOUTCLKFABRIC;
    output RXOUTCLKPCS;
    output RXPHALIGNDONE;
    output RXPHALIGNERR;
    output RXPMARESETDONE;
    output RXPRBSERR;
    output RXPRBSLOCKED;
    output RXPRGDIVRESETDONE;
    output RXRATEDONE;
    output RXRECCLKOUT;
    output RXRESETDONE;
    output RXSLIDERDY;
    output RXSLIPDONE;
    output RXSLIPOUTCLKRDY;
    output RXSLIPPMARDY;
    output [1:0] RXSTARTOFSEQ;
    output [2:0] RXSTATUS;
    output RXSYNCDONE;
    output RXSYNCOUT;
    output RXVALID;
    output [1:0] TXBUFSTATUS;
    output TXCOMFINISH;
    output TXDCCDONE;
    output TXDLYSRESETDONE;
    output TXOUTCLK;
    output TXOUTCLKFABRIC;
    output TXOUTCLKPCS;
    output TXPHALIGNDONE;
    output TXPHINITDONE;
    output TXPMARESETDONE;
    output TXPRGDIVRESETDONE;
    output TXRATEDONE;
    output TXRESETDONE;
    output TXSYNCDONE;
    output TXSYNCOUT;
    input CDRSTEPDIR;
    input CDRSTEPSQ;
    input CDRSTEPSX;
    input CFGRESET;
    input CLKRSVD0;
    input CLKRSVD1;
    input CPLLFREQLOCK;
    input CPLLLOCKDETCLK;
    input CPLLLOCKEN;
    input CPLLPD;
    input [2:0] CPLLREFCLKSEL;
    input CPLLRESET;
    input DMONFIFORESET;
    input DMONITORCLK;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input EYESCANRESET;
    input EYESCANTRIGGER;
    input FREQOS;
    input GTGREFCLK;
    input GTNORTHREFCLK0;
    input GTNORTHREFCLK1;
    input GTREFCLK0;
    input GTREFCLK1;
    input [15:0] GTRSVD;
    input GTRXRESET;
    input GTRXRESETSEL;
    input GTSOUTHREFCLK0;
    input GTSOUTHREFCLK1;
    input GTTXRESET;
    input GTTXRESETSEL;
    input GTYRXN;
    input GTYRXP;
    input INCPCTRL;
    input [2:0] LOOPBACK;
    input PCIEEQRXEQADAPTDONE;
    input PCIERSTIDLE;
    input PCIERSTTXSYNCSTART;
    input PCIEUSERRATEDONE;
    input [15:0] PCSRSVDIN;
    input QPLL0CLK;
    input QPLL0FREQLOCK;
    input QPLL0REFCLK;
    input QPLL1CLK;
    input QPLL1FREQLOCK;
    input QPLL1REFCLK;
    input RESETOVRD;
    input RX8B10BEN;
    input RXAFECFOKEN;
    input RXBUFRESET;
    input RXCDRFREQRESET;
    input RXCDRHOLD;
    input RXCDROVRDEN;
    input RXCDRRESET;
    input RXCHBONDEN;
    input [4:0] RXCHBONDI;
    input [2:0] RXCHBONDLEVEL;
    input RXCHBONDMASTER;
    input RXCHBONDSLAVE;
    input RXCKCALRESET;
    input [6:0] RXCKCALSTART;
    input RXCOMMADETEN;
    input RXDFEAGCHOLD;
    input RXDFEAGCOVRDEN;
    input [3:0] RXDFECFOKFCNUM;
    input RXDFECFOKFEN;
    input RXDFECFOKFPULSE;
    input RXDFECFOKHOLD;
    input RXDFECFOKOVREN;
    input RXDFEKHHOLD;
    input RXDFEKHOVRDEN;
    input RXDFELFHOLD;
    input RXDFELFOVRDEN;
    input RXDFELPMRESET;
    input RXDFETAP10HOLD;
    input RXDFETAP10OVRDEN;
    input RXDFETAP11HOLD;
    input RXDFETAP11OVRDEN;
    input RXDFETAP12HOLD;
    input RXDFETAP12OVRDEN;
    input RXDFETAP13HOLD;
    input RXDFETAP13OVRDEN;
    input RXDFETAP14HOLD;
    input RXDFETAP14OVRDEN;
    input RXDFETAP15HOLD;
    input RXDFETAP15OVRDEN;
    input RXDFETAP2HOLD;
    input RXDFETAP2OVRDEN;
    input RXDFETAP3HOLD;
    input RXDFETAP3OVRDEN;
    input RXDFETAP4HOLD;
    input RXDFETAP4OVRDEN;
    input RXDFETAP5HOLD;
    input RXDFETAP5OVRDEN;
    input RXDFETAP6HOLD;
    input RXDFETAP6OVRDEN;
    input RXDFETAP7HOLD;
    input RXDFETAP7OVRDEN;
    input RXDFETAP8HOLD;
    input RXDFETAP8OVRDEN;
    input RXDFETAP9HOLD;
    input RXDFETAP9OVRDEN;
    input RXDFEUTHOLD;
    input RXDFEUTOVRDEN;
    input RXDFEVPHOLD;
    input RXDFEVPOVRDEN;
    input RXDFEXYDEN;
    input RXDLYBYPASS;
    input RXDLYEN;
    input RXDLYOVRDEN;
    input RXDLYSRESET;
    input [1:0] RXELECIDLEMODE;
    input RXEQTRAINING;
    input RXGEARBOXSLIP;
    input RXLATCLK;
    input RXLPMEN;
    input RXLPMGCHOLD;
    input RXLPMGCOVRDEN;
    input RXLPMHFHOLD;
    input RXLPMHFOVRDEN;
    input RXLPMLFHOLD;
    input RXLPMLFKLOVRDEN;
    input RXLPMOSHOLD;
    input RXLPMOSOVRDEN;
    input RXMCOMMAALIGNEN;
    input [1:0] RXMONITORSEL;
    input RXOOBRESET;
    input RXOSCALRESET;
    input RXOSHOLD;
    input RXOSOVRDEN;
    input [2:0] RXOUTCLKSEL;
    input RXPCOMMAALIGNEN;
    input RXPCSRESET;
    input [1:0] RXPD;
    input RXPHALIGN;
    input RXPHALIGNEN;
    input RXPHDLYPD;
    input RXPHDLYRESET;
    input [1:0] RXPLLCLKSEL;
    input RXPMARESET;
    input RXPOLARITY;
    input RXPRBSCNTRESET;
    input [3:0] RXPRBSSEL;
    input RXPROGDIVRESET;
    input [2:0] RXRATE;
    input RXRATEMODE;
    input RXSLIDE;
    input RXSLIPOUTCLK;
    input RXSLIPPMA;
    input RXSYNCALLIN;
    input RXSYNCIN;
    input RXSYNCMODE;
    input [1:0] RXSYSCLKSEL;
    input RXTERMINATION;
    input RXUSERRDY;
    input RXUSRCLK;
    input RXUSRCLK2;
    input SIGVALIDCLK;
    input [19:0] TSTIN;
    input [7:0] TX8B10BBYPASS;
    input TX8B10BEN;
    input TXCOMINIT;
    input TXCOMSAS;
    input TXCOMWAKE;
    input [15:0] TXCTRL0;
    input [15:0] TXCTRL1;
    input [7:0] TXCTRL2;
    input [127:0] TXDATA;
    input [7:0] TXDATAEXTENDRSVD;
    input TXDCCFORCESTART;
    input TXDCCRESET;
    input [1:0] TXDEEMPH;
    input TXDETECTRX;
    input [4:0] TXDIFFCTRL;
    input TXDLYBYPASS;
    input TXDLYEN;
    input TXDLYHOLD;
    input TXDLYOVRDEN;
    input TXDLYSRESET;
    input TXDLYUPDOWN;
    input TXELECIDLE;
    input [5:0] TXHEADER;
    input TXINHIBIT;
    input TXLATCLK;
    input TXLFPSTRESET;
    input TXLFPSU2LPEXIT;
    input TXLFPSU3WAKE;
    input [6:0] TXMAINCURSOR;
    input [2:0] TXMARGIN;
    input TXMUXDCDEXHOLD;
    input TXMUXDCDORWREN;
    input TXONESZEROS;
    input [2:0] TXOUTCLKSEL;
    input TXPCSRESET;
    input [1:0] TXPD;
    input TXPDELECIDLEMODE;
    input TXPHALIGN;
    input TXPHALIGNEN;
    input TXPHDLYPD;
    input TXPHDLYRESET;
    input TXPHDLYTSTCLK;
    input TXPHINIT;
    input TXPHOVRDEN;
    input TXPIPPMEN;
    input TXPIPPMOVRDEN;
    input TXPIPPMPD;
    input TXPIPPMSEL;
    input [4:0] TXPIPPMSTEPSIZE;
    input TXPISOPD;
    input [1:0] TXPLLCLKSEL;
    input TXPMARESET;
    input TXPOLARITY;
    input [4:0] TXPOSTCURSOR;
    input TXPRBSFORCEERR;
    input [3:0] TXPRBSSEL;
    input [4:0] TXPRECURSOR;
    input TXPROGDIVRESET;
    input [2:0] TXRATE;
    input TXRATEMODE;
    input [6:0] TXSEQUENCE;
    input TXSWING;
    input TXSYNCALLIN;
    input TXSYNCIN;
    input TXSYNCMODE;
    input [1:0] TXSYSCLKSEL;
    input TXUSERRDY;
    input TXUSRCLK;
    input TXUSRCLK2;
endmodule

module GTYE4_COMMON (...);
    parameter [0:0] AEN_QPLL0_FBDIV = 1'b1;
    parameter [0:0] AEN_QPLL1_FBDIV = 1'b1;
    parameter [0:0] AEN_SDM0TOGGLE = 1'b0;
    parameter [0:0] AEN_SDM1TOGGLE = 1'b0;
    parameter [0:0] A_SDM0TOGGLE = 1'b0;
    parameter [8:0] A_SDM1DATA_HIGH = 9'b000000000;
    parameter [15:0] A_SDM1DATA_LOW = 16'b0000000000000000;
    parameter [0:0] A_SDM1TOGGLE = 1'b0;
    parameter [15:0] BIAS_CFG0 = 16'h0000;
    parameter [15:0] BIAS_CFG1 = 16'h0000;
    parameter [15:0] BIAS_CFG2 = 16'h0000;
    parameter [15:0] BIAS_CFG3 = 16'h0000;
    parameter [15:0] BIAS_CFG4 = 16'h0000;
    parameter [15:0] BIAS_CFG_RSVD = 16'h0000;
    parameter [15:0] COMMON_CFG0 = 16'h0000;
    parameter [15:0] COMMON_CFG1 = 16'h0000;
    parameter [15:0] POR_CFG = 16'h0000;
    parameter [15:0] PPF0_CFG = 16'h0F00;
    parameter [15:0] PPF1_CFG = 16'h0F00;
    parameter QPLL0CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL0_CFG0 = 16'h391C;
    parameter [15:0] QPLL0_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL0_CFG2 = 16'h0F80;
    parameter [15:0] QPLL0_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL0_CFG3 = 16'h0120;
    parameter [15:0] QPLL0_CFG4 = 16'h0002;
    parameter [9:0] QPLL0_CP = 10'b0000011111;
    parameter [9:0] QPLL0_CP_G3 = 10'b0000011111;
    parameter integer QPLL0_FBDIV = 66;
    parameter integer QPLL0_FBDIV_G3 = 80;
    parameter [15:0] QPLL0_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL0_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL0_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL0_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL0_LPF = 10'b1011111111;
    parameter [9:0] QPLL0_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL0_PCI_EN = 1'b0;
    parameter [0:0] QPLL0_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL0_REFCLK_DIV = 1;
    parameter [15:0] QPLL0_SDM_CFG0 = 16'h0040;
    parameter [15:0] QPLL0_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL0_SDM_CFG2 = 16'h0000;
    parameter QPLL1CLKOUT_RATE = "FULL";
    parameter [15:0] QPLL1_CFG0 = 16'h691C;
    parameter [15:0] QPLL1_CFG1 = 16'h0020;
    parameter [15:0] QPLL1_CFG1_G3 = 16'h0020;
    parameter [15:0] QPLL1_CFG2 = 16'h0F80;
    parameter [15:0] QPLL1_CFG2_G3 = 16'h0F80;
    parameter [15:0] QPLL1_CFG3 = 16'h0120;
    parameter [15:0] QPLL1_CFG4 = 16'h0002;
    parameter [9:0] QPLL1_CP = 10'b0000011111;
    parameter [9:0] QPLL1_CP_G3 = 10'b0000011111;
    parameter integer QPLL1_FBDIV = 66;
    parameter integer QPLL1_FBDIV_G3 = 80;
    parameter [15:0] QPLL1_INIT_CFG0 = 16'h0000;
    parameter [7:0] QPLL1_INIT_CFG1 = 8'h00;
    parameter [15:0] QPLL1_LOCK_CFG = 16'h01E8;
    parameter [15:0] QPLL1_LOCK_CFG_G3 = 16'h21E8;
    parameter [9:0] QPLL1_LPF = 10'b1011111111;
    parameter [9:0] QPLL1_LPF_G3 = 10'b1111111111;
    parameter [0:0] QPLL1_PCI_EN = 1'b0;
    parameter [0:0] QPLL1_RATE_SW_USE_DRP = 1'b0;
    parameter integer QPLL1_REFCLK_DIV = 1;
    parameter [15:0] QPLL1_SDM_CFG0 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG1 = 16'h0000;
    parameter [15:0] QPLL1_SDM_CFG2 = 16'h0000;
    parameter [15:0] RSVD_ATTR0 = 16'h0000;
    parameter [15:0] RSVD_ATTR1 = 16'h0000;
    parameter [15:0] RSVD_ATTR2 = 16'h0000;
    parameter [15:0] RSVD_ATTR3 = 16'h0000;
    parameter [1:0] RXRECCLKOUT0_SEL = 2'b00;
    parameter [1:0] RXRECCLKOUT1_SEL = 2'b00;
    parameter [0:0] SARC_ENB = 1'b0;
    parameter [0:0] SARC_SEL = 1'b0;
    parameter [15:0] SDM0INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM0INITSEED0_1 = 9'b000000000;
    parameter [15:0] SDM1INITSEED0_0 = 16'b0000000000000000;
    parameter [8:0] SDM1INITSEED0_1 = 9'b000000000;
    parameter SIM_MODE = "FAST";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [15:0] UB_CFG0 = 16'h0000;
    parameter [15:0] UB_CFG1 = 16'h0000;
    parameter [15:0] UB_CFG2 = 16'h0000;
    parameter [15:0] UB_CFG3 = 16'h0000;
    parameter [15:0] UB_CFG4 = 16'h0000;
    parameter [15:0] UB_CFG5 = 16'h0400;
    parameter [15:0] UB_CFG6 = 16'h0000;
    output [15:0] DRPDO;
    output DRPRDY;
    output [7:0] PMARSVDOUT0;
    output [7:0] PMARSVDOUT1;
    output QPLL0FBCLKLOST;
    output QPLL0LOCK;
    output QPLL0OUTCLK;
    output QPLL0OUTREFCLK;
    output QPLL0REFCLKLOST;
    output QPLL1FBCLKLOST;
    output QPLL1LOCK;
    output QPLL1OUTCLK;
    output QPLL1OUTREFCLK;
    output QPLL1REFCLKLOST;
    output [7:0] QPLLDMONITOR0;
    output [7:0] QPLLDMONITOR1;
    output REFCLKOUTMONITOR0;
    output REFCLKOUTMONITOR1;
    output [1:0] RXRECCLK0SEL;
    output [1:0] RXRECCLK1SEL;
    output [3:0] SDM0FINALOUT;
    output [14:0] SDM0TESTDATA;
    output [3:0] SDM1FINALOUT;
    output [14:0] SDM1TESTDATA;
    output [15:0] UBDADDR;
    output UBDEN;
    output [15:0] UBDI;
    output UBDWE;
    output UBMDMTDO;
    output UBRSVDOUT;
    output UBTXUART;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input [15:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input GTGREFCLK0;
    input GTGREFCLK1;
    input GTNORTHREFCLK00;
    input GTNORTHREFCLK01;
    input GTNORTHREFCLK10;
    input GTNORTHREFCLK11;
    input GTREFCLK00;
    input GTREFCLK01;
    input GTREFCLK10;
    input GTREFCLK11;
    input GTSOUTHREFCLK00;
    input GTSOUTHREFCLK01;
    input GTSOUTHREFCLK10;
    input GTSOUTHREFCLK11;
    input [2:0] PCIERATEQPLL0;
    input [2:0] PCIERATEQPLL1;
    input [7:0] PMARSVD0;
    input [7:0] PMARSVD1;
    input QPLL0CLKRSVD0;
    input QPLL0CLKRSVD1;
    input [7:0] QPLL0FBDIV;
    input QPLL0LOCKDETCLK;
    input QPLL0LOCKEN;
    input QPLL0PD;
    input [2:0] QPLL0REFCLKSEL;
    input QPLL0RESET;
    input QPLL1CLKRSVD0;
    input QPLL1CLKRSVD1;
    input [7:0] QPLL1FBDIV;
    input QPLL1LOCKDETCLK;
    input QPLL1LOCKEN;
    input QPLL1PD;
    input [2:0] QPLL1REFCLKSEL;
    input QPLL1RESET;
    input [7:0] QPLLRSVD1;
    input [4:0] QPLLRSVD2;
    input [4:0] QPLLRSVD3;
    input [7:0] QPLLRSVD4;
    input RCALENB;
    input [24:0] SDM0DATA;
    input SDM0RESET;
    input SDM0TOGGLE;
    input [1:0] SDM0WIDTH;
    input [24:0] SDM1DATA;
    input SDM1RESET;
    input SDM1TOGGLE;
    input [1:0] SDM1WIDTH;
    input UBCFGSTREAMEN;
    input [15:0] UBDO;
    input UBDRDY;
    input UBENABLE;
    input [1:0] UBGPI;
    input [1:0] UBINTR;
    input UBIOLMBRST;
    input UBMBRST;
    input UBMDMCAPTURE;
    input UBMDMDBGRST;
    input UBMDMDBGUPDATE;
    input [3:0] UBMDMREGEN;
    input UBMDMSHIFT;
    input UBMDMSYSRST;
    input UBMDMTCK;
    input UBMDMTDI;
endmodule

module IBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [1:0] REFCLK_HROW_CK_SEL = 2'b00;
    parameter [1:0] REFCLK_ICNTL_RX = 2'b00;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module OBUFDS_GTE4 (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTE4_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter [4:0] REFCLK_ICNTL_TX = 5'b00000;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
    input [1:0] RXRECCLK_SEL;
endmodule

module GTM_DUAL (...);
    parameter [15:0] A_CFG = 16'b0000100001000000;
    parameter [15:0] A_SDM_DATA_CFG0 = 16'b0000000011010000;
    parameter [15:0] A_SDM_DATA_CFG1 = 16'b0000000011010000;
    parameter [15:0] BIAS_CFG0 = 16'b0000000000000000;
    parameter [15:0] BIAS_CFG1 = 16'b0000000000000000;
    parameter [15:0] BIAS_CFG2 = 16'b0001000000000000;
    parameter [15:0] BIAS_CFG3 = 16'b0000000000000001;
    parameter [15:0] BIAS_CFG4 = 16'b0000000000000000;
    parameter [15:0] BIAS_CFG5 = 16'b0000000000000000;
    parameter [15:0] BIAS_CFG6 = 16'b0000000010000000;
    parameter [15:0] BIAS_CFG7 = 16'b0000000000000000;
    parameter [15:0] CH0_A_CH_CFG0 = 16'b0000000000000011;
    parameter [15:0] CH0_A_CH_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH0_A_CH_CFG2 = 16'b0111101111110000;
    parameter [15:0] CH0_A_CH_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH0_A_CH_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH0_A_CH_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH0_A_CH_CFG6 = 16'b0000000000000000;
    parameter [15:0] CH0_RST_LP_CFG0 = 16'b0001000000010000;
    parameter [15:0] CH0_RST_LP_CFG1 = 16'b0011001000010000;
    parameter [15:0] CH0_RST_LP_CFG2 = 16'b0110010100000100;
    parameter [15:0] CH0_RST_LP_CFG3 = 16'b0011001000010000;
    parameter [15:0] CH0_RST_LP_CFG4 = 16'b0000000001000100;
    parameter [15:0] CH0_RST_LP_ID_CFG0 = 16'b0011000001110000;
    parameter [15:0] CH0_RST_LP_ID_CFG1 = 16'b0001000000010000;
    parameter [15:0] CH0_RST_TIME_CFG0 = 16'b0000010000100001;
    parameter [15:0] CH0_RST_TIME_CFG1 = 16'b0000010000100001;
    parameter [15:0] CH0_RST_TIME_CFG2 = 16'b0000010000100001;
    parameter [15:0] CH0_RST_TIME_CFG3 = 16'b0000010000100000;
    parameter [15:0] CH0_RST_TIME_CFG4 = 16'b0000010000100001;
    parameter [15:0] CH0_RST_TIME_CFG5 = 16'b0000000000000001;
    parameter [15:0] CH0_RST_TIME_CFG6 = 16'b0000000000100001;
    parameter [15:0] CH0_RX_ADC_CFG0 = 16'b0011010010001111;
    parameter [15:0] CH0_RX_ADC_CFG1 = 16'b0011111001010101;
    parameter [15:0] CH0_RX_ANA_CFG0 = 16'b1000000000011101;
    parameter [15:0] CH0_RX_ANA_CFG1 = 16'b1110100010000000;
    parameter [15:0] CH0_RX_ANA_CFG2 = 16'b0000000010001010;
    parameter [15:0] CH0_RX_APT_CFG0A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG0B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG10A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG10B = 16'b0000000001010000;
    parameter [15:0] CH0_RX_APT_CFG11A = 16'b0000000001000000;
    parameter [15:0] CH0_RX_APT_CFG11B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG12A = 16'b0000000001010000;
    parameter [15:0] CH0_RX_APT_CFG12B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG13A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG13B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG14A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG14B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG15A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG15B = 16'b0000100000000000;
    parameter [15:0] CH0_RX_APT_CFG16A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG16B = 16'b0010000000000000;
    parameter [15:0] CH0_RX_APT_CFG17A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG17B = 16'b0001000001000000;
    parameter [15:0] CH0_RX_APT_CFG18A = 16'b0000100000100000;
    parameter [15:0] CH0_RX_APT_CFG18B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG19A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG19B = 16'b0000100000000000;
    parameter [15:0] CH0_RX_APT_CFG1A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG1B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG20A = 16'b1110000000100000;
    parameter [15:0] CH0_RX_APT_CFG20B = 16'b0000000001000000;
    parameter [15:0] CH0_RX_APT_CFG21A = 16'b0001000000000100;
    parameter [15:0] CH0_RX_APT_CFG21B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG22A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG22B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG23A = 16'b0000100000000000;
    parameter [15:0] CH0_RX_APT_CFG23B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG24A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG24B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG25A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG25B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG26A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG26B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG27A = 16'b0100000000000000;
    parameter [15:0] CH0_RX_APT_CFG27B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG28A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_APT_CFG28B = 16'b1000000000000000;
    parameter [15:0] CH0_RX_APT_CFG2A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG2B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG3A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG3B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG4A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG4B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG5A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG5B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG6A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG6B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG7A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG7B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG8A = 16'b0000100000000000;
    parameter [15:0] CH0_RX_APT_CFG8B = 16'b0000100000000000;
    parameter [15:0] CH0_RX_APT_CFG9A = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CFG9B = 16'b0000000001110000;
    parameter [15:0] CH0_RX_APT_CTRL_CFG2 = 16'b0000000000000100;
    parameter [15:0] CH0_RX_APT_CTRL_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CAL_CFG0A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CAL_CFG0B = 16'b0011001100110000;
    parameter [15:0] CH0_RX_CAL_CFG1A = 16'b1110111011100001;
    parameter [15:0] CH0_RX_CAL_CFG1B = 16'b1111111100000100;
    parameter [15:0] CH0_RX_CAL_CFG2A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CAL_CFG2B = 16'b0011000000000000;
    parameter [15:0] CH0_RX_CDR_CFG0A = 16'b0000000000000011;
    parameter [15:0] CH0_RX_CDR_CFG0B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CDR_CFG1A = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CDR_CFG1B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CDR_CFG2A = 16'b1001000101100100;
    parameter [15:0] CH0_RX_CDR_CFG2B = 16'b0000000100100100;
    parameter [15:0] CH0_RX_CDR_CFG3A = 16'b0101110011110110;
    parameter [15:0] CH0_RX_CDR_CFG3B = 16'b0000000000001011;
    parameter [15:0] CH0_RX_CDR_CFG4A = 16'b0000000000000110;
    parameter [15:0] CH0_RX_CDR_CFG4B = 16'b0000000000000000;
    parameter [15:0] CH0_RX_CLKGN_CFG0 = 16'b1100000000000000;
    parameter [15:0] CH0_RX_CLKGN_CFG1 = 16'b0000000110000000;
    parameter [15:0] CH0_RX_CTLE_CFG0 = 16'b0011010010001000;
    parameter [15:0] CH0_RX_CTLE_CFG1 = 16'b0010000000100010;
    parameter [15:0] CH0_RX_CTLE_CFG2 = 16'b0000101000000000;
    parameter [15:0] CH0_RX_CTLE_CFG3 = 16'b1111001001000000;
    parameter [15:0] CH0_RX_DSP_CFG = 16'b0000000000000000;
    parameter [15:0] CH0_RX_MON_CFG = 16'b0000000000000000;
    parameter [15:0] CH0_RX_PAD_CFG0 = 16'b0001111000000000;
    parameter [15:0] CH0_RX_PAD_CFG1 = 16'b0001100000001010;
    parameter [15:0] CH0_RX_PCS_CFG0 = 16'b0000000100000000;
    parameter [15:0] CH0_RX_PCS_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_ANA_CFG0 = 16'b0000001010101111;
    parameter [15:0] CH0_TX_ANA_CFG1 = 16'b0000000100000000;
    parameter [15:0] CH0_TX_ANA_CFG2 = 16'b1000000000010100;
    parameter [15:0] CH0_TX_ANA_CFG3 = 16'b0000101000100010;
    parameter [15:0] CH0_TX_ANA_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_CAL_CFG0 = 16'b0000000000100000;
    parameter [15:0] CH0_TX_CAL_CFG1 = 16'b0000000001000000;
    parameter [15:0] CH0_TX_DRV_CFG0 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_DRV_CFG1 = 16'b0000000000100111;
    parameter [15:0] CH0_TX_DRV_CFG2 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_DRV_CFG3 = 16'b0110110000000000;
    parameter [15:0] CH0_TX_DRV_CFG4 = 16'b0000000011000101;
    parameter [15:0] CH0_TX_DRV_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_LPBK_CFG0 = 16'b0000000000000011;
    parameter [15:0] CH0_TX_LPBK_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG0 = 16'b0000000101100000;
    parameter [15:0] CH0_TX_PCS_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG10 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG11 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG12 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG13 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG14 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG15 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG16 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG17 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG2 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG6 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG7 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG8 = 16'b0000000000000000;
    parameter [15:0] CH0_TX_PCS_CFG9 = 16'b0000000000000000;
    parameter [15:0] CH1_A_CH_CFG0 = 16'b0000000000000011;
    parameter [15:0] CH1_A_CH_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH1_A_CH_CFG2 = 16'b0111101111110000;
    parameter [15:0] CH1_A_CH_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH1_A_CH_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH1_A_CH_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH1_A_CH_CFG6 = 16'b0000000000000000;
    parameter [15:0] CH1_RST_LP_CFG0 = 16'b0001000000010000;
    parameter [15:0] CH1_RST_LP_CFG1 = 16'b0011001000010000;
    parameter [15:0] CH1_RST_LP_CFG2 = 16'b0110010100000100;
    parameter [15:0] CH1_RST_LP_CFG3 = 16'b0011001000010000;
    parameter [15:0] CH1_RST_LP_CFG4 = 16'b0000000001000100;
    parameter [15:0] CH1_RST_LP_ID_CFG0 = 16'b0011000001110000;
    parameter [15:0] CH1_RST_LP_ID_CFG1 = 16'b0001000000010000;
    parameter [15:0] CH1_RST_TIME_CFG0 = 16'b0000010000100001;
    parameter [15:0] CH1_RST_TIME_CFG1 = 16'b0000010000100001;
    parameter [15:0] CH1_RST_TIME_CFG2 = 16'b0000010000100001;
    parameter [15:0] CH1_RST_TIME_CFG3 = 16'b0000010000100000;
    parameter [15:0] CH1_RST_TIME_CFG4 = 16'b0000010000100001;
    parameter [15:0] CH1_RST_TIME_CFG5 = 16'b0000000000000001;
    parameter [15:0] CH1_RST_TIME_CFG6 = 16'b0000000000100001;
    parameter [15:0] CH1_RX_ADC_CFG0 = 16'b0011010010001111;
    parameter [15:0] CH1_RX_ADC_CFG1 = 16'b0011111001010101;
    parameter [15:0] CH1_RX_ANA_CFG0 = 16'b1000000000011101;
    parameter [15:0] CH1_RX_ANA_CFG1 = 16'b1110100010000000;
    parameter [15:0] CH1_RX_ANA_CFG2 = 16'b0000000010001010;
    parameter [15:0] CH1_RX_APT_CFG0A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG0B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG10A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG10B = 16'b0000000001010000;
    parameter [15:0] CH1_RX_APT_CFG11A = 16'b0000000001000000;
    parameter [15:0] CH1_RX_APT_CFG11B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG12A = 16'b0000000001010000;
    parameter [15:0] CH1_RX_APT_CFG12B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG13A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG13B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG14A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG14B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG15A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG15B = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG16A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG16B = 16'b0010000000000000;
    parameter [15:0] CH1_RX_APT_CFG17A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG17B = 16'b0001000001000000;
    parameter [15:0] CH1_RX_APT_CFG18A = 16'b0000100000100000;
    parameter [15:0] CH1_RX_APT_CFG18B = 16'b0000100010000000;
    parameter [15:0] CH1_RX_APT_CFG19A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG19B = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG1A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG1B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG20A = 16'b1110000000100000;
    parameter [15:0] CH1_RX_APT_CFG20B = 16'b0000000001000000;
    parameter [15:0] CH1_RX_APT_CFG21A = 16'b0001000000000100;
    parameter [15:0] CH1_RX_APT_CFG21B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG22A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG22B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG23A = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG23B = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG24A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG24B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG25A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG25B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG26A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG26B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG27A = 16'b0100000000000000;
    parameter [15:0] CH1_RX_APT_CFG27B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG28A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_APT_CFG28B = 16'b1000000000000000;
    parameter [15:0] CH1_RX_APT_CFG2A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG2B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG3A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG3B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG4A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG4B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG5A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG5B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG6A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG6B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG7A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG7B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG8A = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG8B = 16'b0000100000000000;
    parameter [15:0] CH1_RX_APT_CFG9A = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CFG9B = 16'b0000000001110000;
    parameter [15:0] CH1_RX_APT_CTRL_CFG2 = 16'b0000000000000100;
    parameter [15:0] CH1_RX_APT_CTRL_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CAL_CFG0A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CAL_CFG0B = 16'b0011001100110000;
    parameter [15:0] CH1_RX_CAL_CFG1A = 16'b1110111011100001;
    parameter [15:0] CH1_RX_CAL_CFG1B = 16'b1111111100000100;
    parameter [15:0] CH1_RX_CAL_CFG2A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CAL_CFG2B = 16'b0011000000000000;
    parameter [15:0] CH1_RX_CDR_CFG0A = 16'b0000000000000011;
    parameter [15:0] CH1_RX_CDR_CFG0B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CDR_CFG1A = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CDR_CFG1B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CDR_CFG2A = 16'b1001000101100100;
    parameter [15:0] CH1_RX_CDR_CFG2B = 16'b0000000100100100;
    parameter [15:0] CH1_RX_CDR_CFG3A = 16'b0101110011110110;
    parameter [15:0] CH1_RX_CDR_CFG3B = 16'b0000000000001011;
    parameter [15:0] CH1_RX_CDR_CFG4A = 16'b0000000000000110;
    parameter [15:0] CH1_RX_CDR_CFG4B = 16'b0000000000000000;
    parameter [15:0] CH1_RX_CLKGN_CFG0 = 16'b1100000000000000;
    parameter [15:0] CH1_RX_CLKGN_CFG1 = 16'b0000000110000000;
    parameter [15:0] CH1_RX_CTLE_CFG0 = 16'b0011010010001000;
    parameter [15:0] CH1_RX_CTLE_CFG1 = 16'b0010000000100010;
    parameter [15:0] CH1_RX_CTLE_CFG2 = 16'b0000101000000000;
    parameter [15:0] CH1_RX_CTLE_CFG3 = 16'b1111001001000000;
    parameter [15:0] CH1_RX_DSP_CFG = 16'b0000000000000000;
    parameter [15:0] CH1_RX_MON_CFG = 16'b0000000000000000;
    parameter [15:0] CH1_RX_PAD_CFG0 = 16'b0001111000000000;
    parameter [15:0] CH1_RX_PAD_CFG1 = 16'b0001100000001010;
    parameter [15:0] CH1_RX_PCS_CFG0 = 16'b0000000100000000;
    parameter [15:0] CH1_RX_PCS_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_ANA_CFG0 = 16'b0000001010101111;
    parameter [15:0] CH1_TX_ANA_CFG1 = 16'b0000000100000000;
    parameter [15:0] CH1_TX_ANA_CFG2 = 16'b1000000000010100;
    parameter [15:0] CH1_TX_ANA_CFG3 = 16'b0000101000100010;
    parameter [15:0] CH1_TX_ANA_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_CAL_CFG0 = 16'b0000000000100000;
    parameter [15:0] CH1_TX_CAL_CFG1 = 16'b0000000001000000;
    parameter [15:0] CH1_TX_DRV_CFG0 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_DRV_CFG1 = 16'b0000000000100111;
    parameter [15:0] CH1_TX_DRV_CFG2 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_DRV_CFG3 = 16'b0110110000000000;
    parameter [15:0] CH1_TX_DRV_CFG4 = 16'b0000000011000101;
    parameter [15:0] CH1_TX_DRV_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_LPBK_CFG0 = 16'b0000000000000011;
    parameter [15:0] CH1_TX_LPBK_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG0 = 16'b0000000101100000;
    parameter [15:0] CH1_TX_PCS_CFG1 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG10 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG11 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG12 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG13 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG14 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG15 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG16 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG17 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG2 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG3 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG4 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG5 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG6 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG7 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG8 = 16'b0000000000000000;
    parameter [15:0] CH1_TX_PCS_CFG9 = 16'b0000000000000000;
    parameter real DATARATE = 10.000;
    parameter [15:0] DRPEN_CFG = 16'b0000000000000000;
    parameter [15:0] FEC_CFG0 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG1 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG10 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG11 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG12 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG13 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG14 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG15 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG16 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG17 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG18 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG19 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG2 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG20 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG21 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG22 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG23 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG24 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG25 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG26 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG27 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG3 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG4 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG5 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG6 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG7 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG8 = 16'b0000000000000000;
    parameter [15:0] FEC_CFG9 = 16'b0000000000000000;
    parameter FEC_MODE = "BYPASS";
    parameter real INS_LOSS_NYQ = 20.000;
    parameter integer INTERFACE_WIDTH = 64;
    parameter MODULATION_MODE = "NRZ";
    parameter [15:0] PLL_CFG0 = 16'b0001100111110000;
    parameter [15:0] PLL_CFG1 = 16'b0000111101110000;
    parameter [15:0] PLL_CFG2 = 16'b1000000111101000;
    parameter [15:0] PLL_CFG3 = 16'b0100000000000000;
    parameter [15:0] PLL_CFG4 = 16'b0111111111101010;
    parameter [15:0] PLL_CFG5 = 16'b0100101100111000;
    parameter [15:0] PLL_CFG6 = 16'b0000000000100101;
    parameter [15:0] PLL_CRS_CTRL_CFG0 = 16'b0000101100100000;
    parameter [15:0] PLL_CRS_CTRL_CFG1 = 16'b1100010111010100;
    parameter [0:0] PLL_IPS_PIN_EN = 1'b1;
    parameter integer PLL_IPS_REFCLK_SEL = 0;
    parameter [0:0] RCALSAP_TESTEN = 1'b0;
    parameter [0:0] RCAL_APROBE = 1'b0;
    parameter [15:0] RST_CFG = 16'b0000000000000010;
    parameter [15:0] RST_PLL_CFG0 = 16'b0111011000010100;
    parameter [15:0] SAP_CFG0 = 16'b0000000000000000;
    parameter [15:0] SDM_CFG0 = 16'b0001100001000000;
    parameter [15:0] SDM_CFG1 = 16'b0000000000000000;
    parameter [15:0] SDM_CFG2 = 16'b0000000000000000;
    parameter [15:0] SDM_SEED_CFG0 = 16'b0000000000000000;
    parameter [15:0] SDM_SEED_CFG1 = 16'b0000000000000000;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS_ES1";
    parameter SIM_RESET_SPEEDUP = "TRUE";
    parameter integer TX_AMPLITUDE_SWING = 250;
    output [27:0] CH0_AXISTDATA;
    output CH0_AXISTLAST;
    output CH0_AXISTVALID;
    output [31:0] CH0_DMONITOROUT;
    output CH0_DMONITOROUTCLK;
    output CH0_GTMTXN;
    output CH0_GTMTXP;
    output [15:0] CH0_PCSRSVDOUT;
    output [15:0] CH0_PMARSVDOUT;
    output CH0_RESETEXCEPTION;
    output [2:0] CH0_RXBUFSTATUS;
    output [255:0] CH0_RXDATA;
    output [3:0] CH0_RXDATAFLAGS;
    output CH0_RXDATAISAM;
    output CH0_RXDATASTART;
    output CH0_RXOUTCLK;
    output CH0_RXPMARESETDONE;
    output CH0_RXPRBSERR;
    output CH0_RXPRBSLOCKED;
    output CH0_RXPRGDIVRESETDONE;
    output CH0_RXPROGDIVCLK;
    output CH0_RXRESETDONE;
    output [1:0] CH0_TXBUFSTATUS;
    output CH0_TXOUTCLK;
    output CH0_TXPMARESETDONE;
    output CH0_TXPRGDIVRESETDONE;
    output CH0_TXPROGDIVCLK;
    output CH0_TXRESETDONE;
    output [27:0] CH1_AXISTDATA;
    output CH1_AXISTLAST;
    output CH1_AXISTVALID;
    output [31:0] CH1_DMONITOROUT;
    output CH1_DMONITOROUTCLK;
    output CH1_GTMTXN;
    output CH1_GTMTXP;
    output [15:0] CH1_PCSRSVDOUT;
    output [15:0] CH1_PMARSVDOUT;
    output CH1_RESETEXCEPTION;
    output [2:0] CH1_RXBUFSTATUS;
    output [255:0] CH1_RXDATA;
    output [3:0] CH1_RXDATAFLAGS;
    output CH1_RXDATAISAM;
    output CH1_RXDATASTART;
    output CH1_RXOUTCLK;
    output CH1_RXPMARESETDONE;
    output CH1_RXPRBSERR;
    output CH1_RXPRBSLOCKED;
    output CH1_RXPRGDIVRESETDONE;
    output CH1_RXPROGDIVCLK;
    output CH1_RXRESETDONE;
    output [1:0] CH1_TXBUFSTATUS;
    output CH1_TXOUTCLK;
    output CH1_TXPMARESETDONE;
    output CH1_TXPRGDIVRESETDONE;
    output CH1_TXPROGDIVCLK;
    output CH1_TXRESETDONE;
    output CLKTESTSIG2PAD;
    output DMONITOROUTPLLCLK;
    output [15:0] DRPDO;
    output DRPRDY;
    output FECRX0ALIGNED;
    output FECRX0CORRCWINC;
    output FECRX0CWINC;
    output FECRX0UNCORRCWINC;
    output FECRX1ALIGNED;
    output FECRX1CORRCWINC;
    output FECRX1CWINC;
    output FECRX1UNCORRCWINC;
    output [7:0] FECRXLN0BITERR0TO1INC;
    output [7:0] FECRXLN0BITERR1TO0INC;
    output [14:0] FECRXLN0DLY;
    output [3:0] FECRXLN0ERRCNTINC;
    output [1:0] FECRXLN0MAPPING;
    output [7:0] FECRXLN1BITERR0TO1INC;
    output [7:0] FECRXLN1BITERR1TO0INC;
    output [14:0] FECRXLN1DLY;
    output [3:0] FECRXLN1ERRCNTINC;
    output [1:0] FECRXLN1MAPPING;
    output [7:0] FECRXLN2BITERR0TO1INC;
    output [7:0] FECRXLN2BITERR1TO0INC;
    output [14:0] FECRXLN2DLY;
    output [3:0] FECRXLN2ERRCNTINC;
    output [1:0] FECRXLN2MAPPING;
    output [7:0] FECRXLN3BITERR0TO1INC;
    output [7:0] FECRXLN3BITERR1TO0INC;
    output [14:0] FECRXLN3DLY;
    output [3:0] FECRXLN3ERRCNTINC;
    output [1:0] FECRXLN3MAPPING;
    output FECTRXLN0LOCK;
    output FECTRXLN1LOCK;
    output FECTRXLN2LOCK;
    output FECTRXLN3LOCK;
    output GTPOWERGOOD;
    output PLLFBCLKLOST;
    output PLLLOCK;
    output PLLREFCLKLOST;
    output PLLREFCLKMONITOR;
    output PLLRESETDONE;
    output [15:0] PLLRSVDOUT;
    output RCALCMP;
    output [4:0] RCALOUT;
    output RXRECCLK0;
    output RXRECCLK1;
    input BGBYPASSB;
    input BGMONITORENB;
    input BGPDB;
    input [4:0] BGRCALOVRD;
    input BGRCALOVRDENB;
    input CH0_AXISEN;
    input CH0_AXISRST;
    input CH0_AXISTRDY;
    input CH0_CFGRESET;
    input CH0_DMONFIFORESET;
    input CH0_DMONITORCLK;
    input CH0_GTMRXN;
    input CH0_GTMRXP;
    input CH0_GTRXRESET;
    input CH0_GTTXRESET;
    input [2:0] CH0_LOOPBACK;
    input [15:0] CH0_PCSRSVDIN;
    input [15:0] CH0_PMARSVDIN;
    input CH0_RESETOVRD;
    input CH0_RXADAPTRESET;
    input CH0_RXADCCALRESET;
    input CH0_RXADCCLKGENRESET;
    input CH0_RXBUFRESET;
    input CH0_RXCDRFREQOS;
    input CH0_RXCDRFRRESET;
    input CH0_RXCDRHOLD;
    input CH0_RXCDRINCPCTRL;
    input CH0_RXCDROVRDEN;
    input CH0_RXCDRPHRESET;
    input CH0_RXDFERESET;
    input CH0_RXDSPRESET;
    input CH0_RXEQTRAINING;
    input CH0_RXEYESCANRESET;
    input CH0_RXFECRESET;
    input [2:0] CH0_RXOUTCLKSEL;
    input CH0_RXPCSRESET;
    input [3:0] CH0_RXPCSRESETMASK;
    input CH0_RXPMARESET;
    input [7:0] CH0_RXPMARESETMASK;
    input CH0_RXPOLARITY;
    input CH0_RXPRBSCNTSTOP;
    input CH0_RXPRBSCSCNTRST;
    input [3:0] CH0_RXPRBSPTN;
    input CH0_RXPROGDIVRESET;
    input CH0_RXQPRBSEN;
    input [1:0] CH0_RXRESETMODE;
    input CH0_RXSPCSEQADV;
    input CH0_RXUSRCLK;
    input CH0_RXUSRCLK2;
    input CH0_RXUSRRDY;
    input CH0_RXUSRSTART;
    input CH0_RXUSRSTOP;
    input CH0_TXCKALRESET;
    input [5:0] CH0_TXCTLFIRDAT;
    input [255:0] CH0_TXDATA;
    input CH0_TXDATASTART;
    input [4:0] CH0_TXDRVAMP;
    input [5:0] CH0_TXEMPMAIN;
    input [4:0] CH0_TXEMPPOST;
    input [4:0] CH0_TXEMPPRE;
    input [3:0] CH0_TXEMPPRE2;
    input CH0_TXFECRESET;
    input CH0_TXINHIBIT;
    input CH0_TXMUXDCDEXHOLD;
    input CH0_TXMUXDCDORWREN;
    input [2:0] CH0_TXOUTCLKSEL;
    input CH0_TXPCSRESET;
    input [1:0] CH0_TXPCSRESETMASK;
    input CH0_TXPMARESET;
    input [1:0] CH0_TXPMARESETMASK;
    input CH0_TXPOLARITY;
    input CH0_TXPRBSINERR;
    input [3:0] CH0_TXPRBSPTN;
    input CH0_TXPROGDIVRESET;
    input CH0_TXQPRBSEN;
    input [1:0] CH0_TXRESETMODE;
    input CH0_TXSPCSEQADV;
    input CH0_TXUSRCLK;
    input CH0_TXUSRCLK2;
    input CH0_TXUSRRDY;
    input CH1_AXISEN;
    input CH1_AXISRST;
    input CH1_AXISTRDY;
    input CH1_CFGRESET;
    input CH1_DMONFIFORESET;
    input CH1_DMONITORCLK;
    input CH1_GTMRXN;
    input CH1_GTMRXP;
    input CH1_GTRXRESET;
    input CH1_GTTXRESET;
    input [2:0] CH1_LOOPBACK;
    input [15:0] CH1_PCSRSVDIN;
    input [15:0] CH1_PMARSVDIN;
    input CH1_RESETOVRD;
    input CH1_RXADAPTRESET;
    input CH1_RXADCCALRESET;
    input CH1_RXADCCLKGENRESET;
    input CH1_RXBUFRESET;
    input CH1_RXCDRFREQOS;
    input CH1_RXCDRFRRESET;
    input CH1_RXCDRHOLD;
    input CH1_RXCDRINCPCTRL;
    input CH1_RXCDROVRDEN;
    input CH1_RXCDRPHRESET;
    input CH1_RXDFERESET;
    input CH1_RXDSPRESET;
    input CH1_RXEQTRAINING;
    input CH1_RXEYESCANRESET;
    input CH1_RXFECRESET;
    input [2:0] CH1_RXOUTCLKSEL;
    input CH1_RXPCSRESET;
    input [3:0] CH1_RXPCSRESETMASK;
    input CH1_RXPMARESET;
    input [7:0] CH1_RXPMARESETMASK;
    input CH1_RXPOLARITY;
    input CH1_RXPRBSCNTSTOP;
    input CH1_RXPRBSCSCNTRST;
    input [3:0] CH1_RXPRBSPTN;
    input CH1_RXPROGDIVRESET;
    input CH1_RXQPRBSEN;
    input [1:0] CH1_RXRESETMODE;
    input CH1_RXSPCSEQADV;
    input CH1_RXUSRCLK;
    input CH1_RXUSRCLK2;
    input CH1_RXUSRRDY;
    input CH1_RXUSRSTART;
    input CH1_RXUSRSTOP;
    input CH1_TXCKALRESET;
    input [5:0] CH1_TXCTLFIRDAT;
    input [255:0] CH1_TXDATA;
    input CH1_TXDATASTART;
    input [4:0] CH1_TXDRVAMP;
    input [5:0] CH1_TXEMPMAIN;
    input [4:0] CH1_TXEMPPOST;
    input [4:0] CH1_TXEMPPRE;
    input [3:0] CH1_TXEMPPRE2;
    input CH1_TXFECRESET;
    input CH1_TXINHIBIT;
    input CH1_TXMUXDCDEXHOLD;
    input CH1_TXMUXDCDORWREN;
    input [2:0] CH1_TXOUTCLKSEL;
    input CH1_TXPCSRESET;
    input [1:0] CH1_TXPCSRESETMASK;
    input CH1_TXPMARESET;
    input [1:0] CH1_TXPMARESETMASK;
    input CH1_TXPOLARITY;
    input CH1_TXPRBSINERR;
    input [3:0] CH1_TXPRBSPTN;
    input CH1_TXPROGDIVRESET;
    input CH1_TXQPRBSEN;
    input [1:0] CH1_TXRESETMODE;
    input CH1_TXSPCSEQADV;
    input CH1_TXUSRCLK;
    input CH1_TXUSRCLK2;
    input CH1_TXUSRRDY;
    input [10:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPRST;
    input DRPWE;
    input FECCTRLRX0BITSLIPFS;
    input FECCTRLRX1BITSLIPFS;
    input GTGREFCLK2PLL;
    input GTNORTHREFCLK;
    input GTREFCLK;
    input GTSOUTHREFCLK;
    input [7:0] PLLFBDIV;
    input PLLMONCLK;
    input PLLPD;
    input [2:0] PLLREFCLKSEL;
    input PLLRESET;
    input PLLRESETBYPASSMODE;
    input [1:0] PLLRESETMASK;
    input [15:0] PLLRSVDIN;
    input RCALENB;
    input [25:0] SDMDATA;
    input SDMTOGGLE;
endmodule

module IBUFDS_GTM (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter integer REFCLK_HROW_CK_SEL = 0;
    parameter integer REFCLK_ICNTL_RX = 0;
    output O;
    output ODIV2;
    input CEB;
    (* iopad_external_pin *)
    input I;
    (* iopad_external_pin *)
    input IB;
endmodule

module OBUFDS_GTM (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter integer REFCLK_ICNTL_TX = 0;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input I;
endmodule

module OBUFDS_GTM_ADV (...);
    parameter [0:0] REFCLK_EN_TX_PATH = 1'b0;
    parameter integer REFCLK_ICNTL_TX = 0;
    parameter [1:0] RXRECCLK_SEL = 2'b00;
    (* iopad_external_pin *)
    output O;
    (* iopad_external_pin *)
    output OB;
    input CEB;
    input [3:0] I;
endmodule

module HSDAC (...);
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter integer XPA_CFG0 = 0;
    parameter integer XPA_CFG1 = 0;
    parameter integer XPA_NUM_DACS = 0;
    parameter integer XPA_NUM_DUCS = 0;
    parameter XPA_PLL_USED = "No";
    parameter integer XPA_SAMPLE_RATE_MSPS = 0;
    output CLK_DAC;
    output [15:0] DOUT;
    output DRDY;
    output PLL_DMON_OUT;
    output PLL_REFCLK_OUT;
    output [15:0] STATUS_COMMON;
    output [15:0] STATUS_DAC0;
    output [15:0] STATUS_DAC1;
    output [15:0] STATUS_DAC2;
    output [15:0] STATUS_DAC3;
    output SYSREF_OUT_NORTH;
    output SYSREF_OUT_SOUTH;
    output VOUT0_N;
    output VOUT0_P;
    output VOUT1_N;
    output VOUT1_P;
    output VOUT2_N;
    output VOUT2_P;
    output VOUT3_N;
    output VOUT3_P;
    input CLK_FIFO_LM;
    input [15:0] CONTROL_COMMON;
    input [15:0] CONTROL_DAC0;
    input [15:0] CONTROL_DAC1;
    input [15:0] CONTROL_DAC2;
    input [15:0] CONTROL_DAC3;
    input DAC_CLK_N;
    input DAC_CLK_P;
    input [11:0] DADDR;
    input [255:0] DATA_DAC0;
    input [255:0] DATA_DAC1;
    input [255:0] DATA_DAC2;
    input [255:0] DATA_DAC3;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input FABRIC_CLK;
    input PLL_MONCLK;
    input PLL_REFCLK_IN;
    input SYSREF_IN_NORTH;
    input SYSREF_IN_SOUTH;
    input SYSREF_N;
    input SYSREF_P;
endmodule

module HSADC (...);
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter integer XPA_CFG0 = 0;
    parameter integer XPA_CFG1 = 0;
    parameter XPA_NUM_ADCS = "0";
    parameter integer XPA_NUM_DDCS = 0;
    parameter XPA_PLL_USED = "No";
    parameter integer XPA_SAMPLE_RATE_MSPS = 0;
    output CLK_ADC;
    output [127:0] DATA_ADC0;
    output [127:0] DATA_ADC1;
    output [127:0] DATA_ADC2;
    output [127:0] DATA_ADC3;
    output [15:0] DOUT;
    output DRDY;
    output PLL_DMON_OUT;
    output PLL_REFCLK_OUT;
    output [15:0] STATUS_ADC0;
    output [15:0] STATUS_ADC1;
    output [15:0] STATUS_ADC2;
    output [15:0] STATUS_ADC3;
    output [15:0] STATUS_COMMON;
    output SYSREF_OUT_NORTH;
    output SYSREF_OUT_SOUTH;
    input ADC_CLK_N;
    input ADC_CLK_P;
    input CLK_FIFO_LM;
    input [15:0] CONTROL_ADC0;
    input [15:0] CONTROL_ADC1;
    input [15:0] CONTROL_ADC2;
    input [15:0] CONTROL_ADC3;
    input [15:0] CONTROL_COMMON;
    input [11:0] DADDR;
    input DCLK;
    input DEN;
    input [15:0] DI;
    input DWE;
    input FABRIC_CLK;
    input PLL_MONCLK;
    input PLL_REFCLK_IN;
    input SYSREF_IN_NORTH;
    input SYSREF_IN_SOUTH;
    input SYSREF_N;
    input SYSREF_P;
    input VIN0_N;
    input VIN0_P;
    input VIN1_N;
    input VIN1_P;
    input VIN2_N;
    input VIN2_P;
    input VIN3_N;
    input VIN3_P;
    input VIN_I01_N;
    input VIN_I01_P;
    input VIN_I23_N;
    input VIN_I23_P;
endmodule

module PCIE_2_1 (...);
    parameter [11:0] AER_BASE_PTR = 12'h140;
    parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [15:0] AER_CAP_ID = 16'h0001;
    parameter AER_CAP_MULTIHEADER = "FALSE";
    parameter [11:0] AER_CAP_NEXTPTR = 12'h178;
    parameter AER_CAP_ON = "FALSE";
    parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000;
    parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
    parameter [3:0] AER_CAP_VERSION = 4'h2;
    parameter ALLOW_X8_GEN2 = "FALSE";
    parameter [31:0] BAR0 = 32'hFFFFFF00;
    parameter [31:0] BAR1 = 32'hFFFF0000;
    parameter [31:0] BAR2 = 32'hFFFF000C;
    parameter [31:0] BAR3 = 32'hFFFFFFFF;
    parameter [31:0] BAR4 = 32'h00000000;
    parameter [31:0] BAR5 = 32'h00000000;
    parameter [7:0] CAPABILITIES_PTR = 8'h40;
    parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
    parameter integer CFG_ECRC_ERR_CPLSTAT = 0;
    parameter [23:0] CLASS_CODE = 24'h000000;
    parameter CMD_INTX_IMPLEMENTED = "TRUE";
    parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
    parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
    parameter [6:0] CRM_MODULE_RSTS = 7'h00;
    parameter DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE";
    parameter DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE";
    parameter DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE";
    parameter DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE";
    parameter DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE";
    parameter [1:0] DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0;
    parameter DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE";
    parameter [1:0] DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0;
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
    parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
    parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
    parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
    parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
    parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
    parameter integer DEV_CAP_RSVD_14_12 = 0;
    parameter integer DEV_CAP_RSVD_17_16 = 0;
    parameter integer DEV_CAP_RSVD_31_29 = 0;
    parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
    parameter DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE";
    parameter DISABLE_ASPM_L1_TIMER = "FALSE";
    parameter DISABLE_BAR_FILTERING = "FALSE";
    parameter DISABLE_ERR_MSG = "FALSE";
    parameter DISABLE_ID_CHECK = "FALSE";
    parameter DISABLE_LANE_REVERSAL = "FALSE";
    parameter DISABLE_LOCKED_FILTER = "FALSE";
    parameter DISABLE_PPM_FILTER = "FALSE";
    parameter DISABLE_RX_POISONED_RESP = "FALSE";
    parameter DISABLE_RX_TC_FILTER = "FALSE";
    parameter DISABLE_SCRAMBLING = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [11:0] DSN_BASE_PTR = 12'h100;
    parameter [15:0] DSN_CAP_ID = 16'h0003;
    parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C;
    parameter DSN_CAP_ON = "TRUE";
    parameter [3:0] DSN_CAP_VERSION = 4'h1;
    parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
    parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
    parameter ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE";
    parameter ENTER_RVRY_EI_L0 = "TRUE";
    parameter EXIT_LOOPBACK_ON_EI = "TRUE";
    parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
    parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
    parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
    parameter [7:0] HEADER_TYPE = 8'h00;
    parameter [4:0] INFER_EI = 5'h00;
    parameter [7:0] INTERRUPT_PIN = 8'h01;
    parameter INTERRUPT_STAT_AUTO = "TRUE";
    parameter IS_SWITCH = "FALSE";
    parameter [9:0] LAST_CONFIG_DWORD = 10'h3FF;
    parameter LINK_CAP_ASPM_OPTIONALITY = "TRUE";
    parameter integer LINK_CAP_ASPM_SUPPORT = 1;
    parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
    parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
    parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
    parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
    parameter integer LINK_CAP_RSVD_23 = 0;
    parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
    parameter integer LINK_CONTROL_RCB = 0;
    parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
    parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
    parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
    parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
    parameter MPS_FORCE = "FALSE";
    parameter [7:0] MSIX_BASE_PTR = 8'h9C;
    parameter [7:0] MSIX_CAP_ID = 8'h11;
    parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
    parameter MSIX_CAP_ON = "FALSE";
    parameter integer MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] MSI_BASE_PTR = 8'h48;
    parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
    parameter [7:0] MSI_CAP_ID = 8'h05;
    parameter integer MSI_CAP_MULTIMSGCAP = 0;
    parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
    parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
    parameter MSI_CAP_ON = "FALSE";
    parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
    parameter integer N_FTS_COMCLK_GEN1 = 255;
    parameter integer N_FTS_COMCLK_GEN2 = 255;
    parameter integer N_FTS_GEN1 = 255;
    parameter integer N_FTS_GEN2 = 255;
    parameter [7:0] PCIE_BASE_PTR = 8'h60;
    parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
    parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
    parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
    parameter [7:0] PCIE_CAP_NEXTPTR = 8'h9C;
    parameter PCIE_CAP_ON = "TRUE";
    parameter integer PCIE_CAP_RSVD_15_14 = 0;
    parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
    parameter integer PCIE_REVISION = 2;
    parameter integer PL_AUTO_CONFIG = 0;
    parameter PL_FAST_TRAIN = "FALSE";
    parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000;
    parameter PM_ASPML0S_TIMEOUT_EN = "FALSE";
    parameter integer PM_ASPML0S_TIMEOUT_FUNC = 0;
    parameter PM_ASPM_FASTEXIT = "FALSE";
    parameter [7:0] PM_BASE_PTR = 8'h40;
    parameter integer PM_CAP_AUXCURRENT = 0;
    parameter PM_CAP_D1SUPPORT = "TRUE";
    parameter PM_CAP_D2SUPPORT = "TRUE";
    parameter PM_CAP_DSI = "FALSE";
    parameter [7:0] PM_CAP_ID = 8'h01;
    parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
    parameter PM_CAP_ON = "TRUE";
    parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
    parameter PM_CAP_PME_CLOCK = "FALSE";
    parameter integer PM_CAP_RSVD_04 = 0;
    parameter integer PM_CAP_VERSION = 3;
    parameter PM_CSR_B2B3 = "FALSE";
    parameter PM_CSR_BPCCEN = "FALSE";
    parameter PM_CSR_NOSOFTRST = "TRUE";
    parameter [7:0] PM_DATA0 = 8'h01;
    parameter [7:0] PM_DATA1 = 8'h01;
    parameter [7:0] PM_DATA2 = 8'h01;
    parameter [7:0] PM_DATA3 = 8'h01;
    parameter [7:0] PM_DATA4 = 8'h01;
    parameter [7:0] PM_DATA5 = 8'h01;
    parameter [7:0] PM_DATA6 = 8'h01;
    parameter [7:0] PM_DATA7 = 8'h01;
    parameter [1:0] PM_DATA_SCALE0 = 2'h1;
    parameter [1:0] PM_DATA_SCALE1 = 2'h1;
    parameter [1:0] PM_DATA_SCALE2 = 2'h1;
    parameter [1:0] PM_DATA_SCALE3 = 2'h1;
    parameter [1:0] PM_DATA_SCALE4 = 2'h1;
    parameter [1:0] PM_DATA_SCALE5 = 2'h1;
    parameter [1:0] PM_DATA_SCALE6 = 2'h1;
    parameter [1:0] PM_DATA_SCALE7 = 2'h1;
    parameter PM_MF = "FALSE";
    parameter [11:0] RBAR_BASE_PTR = 12'h178;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00;
    parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00;
    parameter [15:0] RBAR_CAP_ID = 16'h0015;
    parameter [2:0] RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX2 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX3 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX4 = 3'h0;
    parameter [2:0] RBAR_CAP_INDEX5 = 3'h0;
    parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000;
    parameter RBAR_CAP_ON = "FALSE";
    parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000;
    parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000;
    parameter [3:0] RBAR_CAP_VERSION = 4'h1;
    parameter [2:0] RBAR_NUM = 3'h1;
    parameter integer RECRC_CHK = 0;
    parameter RECRC_CHK_TRIM = "FALSE";
    parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
    parameter [1:0] RP_AUTO_SPD = 2'h1;
    parameter [4:0] RP_AUTO_SPD_LOOPCNT = 5'h1F;
    parameter SELECT_DLL_IF = "FALSE";
    parameter SIM_VERSION = "1.0";
    parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
    parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
    parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
    parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
    parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
    parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
    parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
    parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
    parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
    parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
    parameter integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
    parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SSL_MESSAGE_AUTO = "FALSE";
    parameter TECRC_EP_INV = "FALSE";
    parameter TL_RBYPASS = "FALSE";
    parameter integer TL_RX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
    parameter TL_TFC_DISABLE = "FALSE";
    parameter TL_TX_CHECKS_DISABLE = "FALSE";
    parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
    parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
    parameter integer TL_TX_RAM_WRITE_LATENCY = 0;
    parameter TRN_DW = "FALSE";
    parameter TRN_NP_FC = "FALSE";
    parameter UPCONFIG_CAPABLE = "TRUE";
    parameter UPSTREAM_FACING = "TRUE";
    parameter UR_ATOMIC = "TRUE";
    parameter UR_CFG1 = "TRUE";
    parameter UR_INV_REQ = "TRUE";
    parameter UR_PRS_RESPONSE = "TRUE";
    parameter USER_CLK2_DIV2 = "FALSE";
    parameter integer USER_CLK_FREQ = 3;
    parameter USE_RID_PINS = "FALSE";
    parameter VC0_CPL_INFINITE = "TRUE";
    parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
    parameter integer VC0_TOTAL_CREDITS_CD = 127;
    parameter integer VC0_TOTAL_CREDITS_CH = 31;
    parameter integer VC0_TOTAL_CREDITS_NPD = 24;
    parameter integer VC0_TOTAL_CREDITS_NPH = 12;
    parameter integer VC0_TOTAL_CREDITS_PD = 288;
    parameter integer VC0_TOTAL_CREDITS_PH = 32;
    parameter integer VC0_TX_LASTPACKET = 31;
    parameter [11:0] VC_BASE_PTR = 12'h10C;
    parameter [15:0] VC_CAP_ID = 16'h0002;
    parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
    parameter VC_CAP_ON = "FALSE";
    parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
    parameter [3:0] VC_CAP_VERSION = 4'h1;
    parameter [11:0] VSEC_BASE_PTR = 12'h128;
    parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
    parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
    parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
    parameter [15:0] VSEC_CAP_ID = 16'h000B;
    parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
    parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140;
    parameter VSEC_CAP_ON = "FALSE";
    parameter [3:0] VSEC_CAP_VERSION = 4'h1;
    output CFGAERECRCCHECKEN;
    output CFGAERECRCGENEN;
    output CFGAERROOTERRCORRERRRECEIVED;
    output CFGAERROOTERRCORRERRREPORTINGEN;
    output CFGAERROOTERRFATALERRRECEIVED;
    output CFGAERROOTERRFATALERRREPORTINGEN;
    output CFGAERROOTERRNONFATALERRRECEIVED;
    output CFGAERROOTERRNONFATALERRREPORTINGEN;
    output CFGBRIDGESERREN;
    output CFGCOMMANDBUSMASTERENABLE;
    output CFGCOMMANDINTERRUPTDISABLE;
    output CFGCOMMANDIOENABLE;
    output CFGCOMMANDMEMENABLE;
    output CFGCOMMANDSERREN;
    output CFGDEVCONTROL2ARIFORWARDEN;
    output CFGDEVCONTROL2ATOMICEGRESSBLOCK;
    output CFGDEVCONTROL2ATOMICREQUESTEREN;
    output CFGDEVCONTROL2CPLTIMEOUTDIS;
    output CFGDEVCONTROL2IDOCPLEN;
    output CFGDEVCONTROL2IDOREQEN;
    output CFGDEVCONTROL2LTREN;
    output CFGDEVCONTROL2TLPPREFIXBLOCK;
    output CFGDEVCONTROLAUXPOWEREN;
    output CFGDEVCONTROLCORRERRREPORTINGEN;
    output CFGDEVCONTROLENABLERO;
    output CFGDEVCONTROLEXTTAGEN;
    output CFGDEVCONTROLFATALERRREPORTINGEN;
    output CFGDEVCONTROLNONFATALREPORTINGEN;
    output CFGDEVCONTROLNOSNOOPEN;
    output CFGDEVCONTROLPHANTOMEN;
    output CFGDEVCONTROLURERRREPORTINGEN;
    output CFGDEVSTATUSCORRERRDETECTED;
    output CFGDEVSTATUSFATALERRDETECTED;
    output CFGDEVSTATUSNONFATALERRDETECTED;
    output CFGDEVSTATUSURDETECTED;
    output CFGERRAERHEADERLOGSETN;
    output CFGERRCPLRDYN;
    output CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFM;
    output CFGINTERRUPTRDYN;
    output CFGLINKCONTROLAUTOBANDWIDTHINTEN;
    output CFGLINKCONTROLBANDWIDTHINTEN;
    output CFGLINKCONTROLCLOCKPMEN;
    output CFGLINKCONTROLCOMMONCLOCK;
    output CFGLINKCONTROLEXTENDEDSYNC;
    output CFGLINKCONTROLHWAUTOWIDTHDIS;
    output CFGLINKCONTROLLINKDISABLE;
    output CFGLINKCONTROLRCB;
    output CFGLINKCONTROLRETRAINLINK;
    output CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
    output CFGLINKSTATUSBANDWIDTHSTATUS;
    output CFGLINKSTATUSDLLACTIVE;
    output CFGLINKSTATUSLINKTRAINING;
    output CFGMGMTRDWRDONEN;
    output CFGMSGRECEIVED;
    output CFGMSGRECEIVEDASSERTINTA;
    output CFGMSGRECEIVEDASSERTINTB;
    output CFGMSGRECEIVEDASSERTINTC;
    output CFGMSGRECEIVEDASSERTINTD;
    output CFGMSGRECEIVEDDEASSERTINTA;
    output CFGMSGRECEIVEDDEASSERTINTB;
    output CFGMSGRECEIVEDDEASSERTINTC;
    output CFGMSGRECEIVEDDEASSERTINTD;
    output CFGMSGRECEIVEDERRCOR;
    output CFGMSGRECEIVEDERRFATAL;
    output CFGMSGRECEIVEDERRNONFATAL;
    output CFGMSGRECEIVEDPMASNAK;
    output CFGMSGRECEIVEDPMETO;
    output CFGMSGRECEIVEDPMETOACK;
    output CFGMSGRECEIVEDPMPME;
    output CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
    output CFGMSGRECEIVEDUNLOCK;
    output CFGPMCSRPMEEN;
    output CFGPMCSRPMESTATUS;
    output CFGPMRCVASREQL1N;
    output CFGPMRCVENTERL1N;
    output CFGPMRCVENTERL23N;
    output CFGPMRCVREQACKN;
    output CFGROOTCONTROLPMEINTEN;
    output CFGROOTCONTROLSYSERRCORRERREN;
    output CFGROOTCONTROLSYSERRFATALERREN;
    output CFGROOTCONTROLSYSERRNONFATALERREN;
    output CFGSLOTCONTROLELECTROMECHILCTLPULSE;
    output CFGTRANSACTION;
    output CFGTRANSACTIONTYPE;
    output DBGSCLRA;
    output DBGSCLRB;
    output DBGSCLRC;
    output DBGSCLRD;
    output DBGSCLRE;
    output DBGSCLRF;
    output DBGSCLRG;
    output DBGSCLRH;
    output DBGSCLRI;
    output DBGSCLRJ;
    output DBGSCLRK;
    output DRPRDY;
    output LL2BADDLLPERR;
    output LL2BADTLPERR;
    output LL2PROTOCOLERR;
    output LL2RECEIVERERR;
    output LL2REPLAYROERR;
    output LL2REPLAYTOERR;
    output LL2SUSPENDOK;
    output LL2TFCINIT1SEQ;
    output LL2TFCINIT2SEQ;
    output LL2TXIDLE;
    output LNKCLKEN;
    output MIMRXREN;
    output MIMRXWEN;
    output MIMTXREN;
    output MIMTXWEN;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0ELECIDLE;
    output PIPETX1COMPLIANCE;
    output PIPETX1ELECIDLE;
    output PIPETX2COMPLIANCE;
    output PIPETX2ELECIDLE;
    output PIPETX3COMPLIANCE;
    output PIPETX3ELECIDLE;
    output PIPETX4COMPLIANCE;
    output PIPETX4ELECIDLE;
    output PIPETX5COMPLIANCE;
    output PIPETX5ELECIDLE;
    output PIPETX6COMPLIANCE;
    output PIPETX6ELECIDLE;
    output PIPETX7COMPLIANCE;
    output PIPETX7ELECIDLE;
    output PIPETXDEEMPH;
    output PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PL2L0REQ;
    output PL2LINKUP;
    output PL2RECEIVERERR;
    output PL2RECOVERY;
    output PL2RXELECIDLE;
    output PL2SUSPENDOK;
    output PLDIRECTEDCHANGEDONE;
    output PLLINKGEN2CAP;
    output PLLINKPARTNERGEN2SUPPORTED;
    output PLLINKUPCFGCAP;
    output PLPHYLNKUPN;
    output PLRECEIVEDHOTRST;
    output PLSELLNKRATE;
    output RECEIVEDFUNCLVLRSTN;
    output TL2ASPMSUSPENDCREDITCHECKOK;
    output TL2ASPMSUSPENDREQ;
    output TL2ERRFCPE;
    output TL2ERRMALFORMED;
    output TL2ERRRXOVERFLOW;
    output TL2PPMSUSPENDOK;
    output TRNLNKUP;
    output TRNRECRCERR;
    output TRNREOF;
    output TRNRERRFWD;
    output TRNRSOF;
    output TRNRSRCDSC;
    output TRNRSRCRDY;
    output TRNTCFGREQ;
    output TRNTDLLPDSTRDY;
    output TRNTERRDROP;
    output USERRSTN;
    output [11:0] DBGVECC;
    output [11:0] PLDBGVEC;
    output [11:0] TRNFCCPLD;
    output [11:0] TRNFCNPD;
    output [11:0] TRNFCPD;
    output [127:0] TRNRD;
    output [12:0] MIMRXRADDR;
    output [12:0] MIMRXWADDR;
    output [12:0] MIMTXRADDR;
    output [12:0] MIMTXWADDR;
    output [15:0] CFGMSGDATA;
    output [15:0] DRPDO;
    output [15:0] PIPETX0DATA;
    output [15:0] PIPETX1DATA;
    output [15:0] PIPETX2DATA;
    output [15:0] PIPETX3DATA;
    output [15:0] PIPETX4DATA;
    output [15:0] PIPETX5DATA;
    output [15:0] PIPETX6DATA;
    output [15:0] PIPETX7DATA;
    output [1:0] CFGLINKCONTROLASPMCONTROL;
    output [1:0] CFGLINKSTATUSCURRENTSPEED;
    output [1:0] CFGPMCSRPOWERSTATE;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PL2RXPMSTATE;
    output [1:0] PLLANEREVERSALMODE;
    output [1:0] PLRXPMSTATE;
    output [1:0] PLSELLNKWIDTH;
    output [1:0] TRNRDLLPSRCRDY;
    output [1:0] TRNRREM;
    output [2:0] CFGDEVCONTROLMAXPAYLOAD;
    output [2:0] CFGDEVCONTROLMAXREADREQ;
    output [2:0] CFGINTERRUPTMMENABLE;
    output [2:0] CFGPCIELINKSTATE;
    output [2:0] PIPETXMARGIN;
    output [2:0] PLINITIALLINKWIDTH;
    output [2:0] PLTXPMSTATE;
    output [31:0] CFGMGMTDO;
    output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL;
    output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH;
    output [3:0] TRNTDSTRDY;
    output [4:0] LL2LINKSTATUS;
    output [5:0] PLLTSSMSTATE;
    output [5:0] TRNTBUFAV;
    output [63:0] DBGVECA;
    output [63:0] DBGVECB;
    output [63:0] TL2ERRHDR;
    output [63:0] TRNRDLLPDATA;
    output [67:0] MIMRXWDATA;
    output [68:0] MIMTXWDATA;
    output [6:0] CFGTRANSACTIONADDR;
    output [6:0] CFGVCTCVCMAP;
    output [7:0] CFGINTERRUPTDO;
    output [7:0] TRNFCCPLH;
    output [7:0] TRNFCNPH;
    output [7:0] TRNFCPH;
    output [7:0] TRNRBARHIT;
    input CFGERRACSN;
    input CFGERRATOMICEGRESSBLOCKEDN;
    input CFGERRCORN;
    input CFGERRCPLABORTN;
    input CFGERRCPLTIMEOUTN;
    input CFGERRCPLUNEXPECTN;
    input CFGERRECRCN;
    input CFGERRINTERNALCORN;
    input CFGERRINTERNALUNCORN;
    input CFGERRLOCKEDN;
    input CFGERRMALFORMEDN;
    input CFGERRMCBLOCKEDN;
    input CFGERRNORECOVERYN;
    input CFGERRPOISONEDN;
    input CFGERRPOSTEDN;
    input CFGERRURN;
    input CFGFORCECOMMONCLOCKOFF;
    input CFGFORCEEXTENDEDSYNCON;
    input CFGINTERRUPTASSERTN;
    input CFGINTERRUPTN;
    input CFGINTERRUPTSTATN;
    input CFGMGMTRDENN;
    input CFGMGMTWRENN;
    input CFGMGMTWRREADONLYN;
    input CFGMGMTWRRW1CASRWN;
    input CFGPMFORCESTATEENN;
    input CFGPMHALTASPML0SN;
    input CFGPMHALTASPML1N;
    input CFGPMSENDPMETON;
    input CFGPMTURNOFFOKN;
    input CFGPMWAKEN;
    input CFGTRNPENDINGN;
    input CMRSTN;
    input CMSTICKYRSTN;
    input DBGSUBMODE;
    input DLRSTN;
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input FUNCLVLRSTN;
    input LL2SENDASREQL1;
    input LL2SENDENTERL1;
    input LL2SENDENTERL23;
    input LL2SENDPMACK;
    input LL2SUSPENDNOW;
    input LL2TLPRCV;
    input PIPECLK;
    input PIPERX0CHANISALIGNED;
    input PIPERX0ELECIDLE;
    input PIPERX0PHYSTATUS;
    input PIPERX0VALID;
    input PIPERX1CHANISALIGNED;
    input PIPERX1ELECIDLE;
    input PIPERX1PHYSTATUS;
    input PIPERX1VALID;
    input PIPERX2CHANISALIGNED;
    input PIPERX2ELECIDLE;
    input PIPERX2PHYSTATUS;
    input PIPERX2VALID;
    input PIPERX3CHANISALIGNED;
    input PIPERX3ELECIDLE;
    input PIPERX3PHYSTATUS;
    input PIPERX3VALID;
    input PIPERX4CHANISALIGNED;
    input PIPERX4ELECIDLE;
    input PIPERX4PHYSTATUS;
    input PIPERX4VALID;
    input PIPERX5CHANISALIGNED;
    input PIPERX5ELECIDLE;
    input PIPERX5PHYSTATUS;
    input PIPERX5VALID;
    input PIPERX6CHANISALIGNED;
    input PIPERX6ELECIDLE;
    input PIPERX6PHYSTATUS;
    input PIPERX6VALID;
    input PIPERX7CHANISALIGNED;
    input PIPERX7ELECIDLE;
    input PIPERX7PHYSTATUS;
    input PIPERX7VALID;
    input PLDIRECTEDLINKAUTON;
    input PLDIRECTEDLINKSPEED;
    input PLDIRECTEDLTSSMNEWVLD;
    input PLDIRECTEDLTSSMSTALL;
    input PLDOWNSTREAMDEEMPHSOURCE;
    input PLRSTN;
    input PLTRANSMITHOTRST;
    input PLUPSTREAMPREFERDEEMPH;
    input SYSRSTN;
    input TL2ASPMSUSPENDCREDITCHECK;
    input TL2PPMSUSPENDREQ;
    input TLRSTN;
    input TRNRDSTRDY;
    input TRNRFCPRET;
    input TRNRNPOK;
    input TRNRNPREQ;
    input TRNTCFGGNT;
    input TRNTDLLPSRCRDY;
    input TRNTECRCGEN;
    input TRNTEOF;
    input TRNTERRFWD;
    input TRNTSOF;
    input TRNTSRCDSC;
    input TRNTSRCRDY;
    input TRNTSTR;
    input USERCLK2;
    input USERCLK;
    input [127:0] CFGERRAERHEADERLOG;
    input [127:0] TRNTD;
    input [15:0] CFGDEVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [15:0] CFGVENDID;
    input [15:0] DRPDI;
    input [15:0] PIPERX0DATA;
    input [15:0] PIPERX1DATA;
    input [15:0] PIPERX2DATA;
    input [15:0] PIPERX3DATA;
    input [15:0] PIPERX4DATA;
    input [15:0] PIPERX5DATA;
    input [15:0] PIPERX6DATA;
    input [15:0] PIPERX7DATA;
    input [1:0] CFGPMFORCESTATE;
    input [1:0] DBGMODE;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PLDIRECTEDLINKCHANGE;
    input [1:0] PLDIRECTEDLINKWIDTH;
    input [1:0] TRNTREM;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] CFGFORCEMPS;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [2:0] PLDBGMODE;
    input [2:0] TRNFCSEL;
    input [31:0] CFGMGMTDI;
    input [31:0] TRNTDLLPDATA;
    input [3:0] CFGMGMTBYTEENN;
    input [47:0] CFGERRTLPCPLHEADER;
    input [4:0] CFGAERINTERRUPTMSGNUM;
    input [4:0] CFGDSDEVICENUMBER;
    input [4:0] CFGPCIECAPINTERRUPTMSGNUM;
    input [4:0] PL2DIRECTEDLSTATE;
    input [5:0] PLDIRECTEDLTSSMNEW;
    input [63:0] CFGDSN;
    input [67:0] MIMRXRDATA;
    input [68:0] MIMTXRDATA;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGINTERRUPTDI;
    input [7:0] CFGPORTNUMBER;
    input [7:0] CFGREVID;
    input [8:0] DRPADDR;
    input [9:0] CFGMGMTDWADDR;
endmodule

module PCIE_3_0 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
    parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [1:0] GEN3_PCS_AUTO_REALIGN = 2'h1;
    parameter GEN3_PCS_RX_ELECIDLE_INTERNAL = "TRUE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [4:0] PF0_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_BIST_REGISTER = 8'h00;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter [15:0] PF0_DEVICE_ID = 16'h0000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
    parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF0_PB_CAP_VER = 4'h1;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter PF0_RBAR_CAP_ENABLE = "FALSE";
    parameter [2:0] PF0_RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] PF0_RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] PF0_RBAR_CAP_INDEX2 = 3'h0;
    parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF0_RBAR_NUM = 3'h1;
    parameter [7:0] PF0_REVISION_ID = 8'h00;
    parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [4:0] PF1_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_BIST_REGISTER = 8'h00;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [15:0] PF1_DEVICE_ID = 16'h0000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
    parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF1_PB_CAP_VER = 4'h1;
    parameter [7:0] PF1_PM_CAP_ID = 8'h01;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
    parameter PF1_RBAR_CAP_ENABLE = "FALSE";
    parameter [2:0] PF1_RBAR_CAP_INDEX0 = 3'h0;
    parameter [2:0] PF1_RBAR_CAP_INDEX1 = 3'h0;
    parameter [2:0] PF1_RBAR_CAP_INDEX2 = 3'h0;
    parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF1_RBAR_NUM = 3'h1;
    parameter [7:0] PF1_REVISION_ID = 8'h00;
    parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
    parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF1_TPHR_CAP_ENABLE = "FALSE";
    parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_SCRAMBLING = "FALSE";
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
    parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
    parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
    parameter integer PL_N_FTS_GEN1 = 255;
    parameter integer PL_N_FTS_GEN2 = 255;
    parameter integer PL_N_FTS_GEN3 = 255;
    parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
    parameter SIM_VERSION = "1.0";
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SRIOV_CAP_ENABLE = "FALSE";
    parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h0000000;
    parameter [11:0] TL_CREDITS_CD = 12'h3E0;
    parameter [7:0] TL_CREDITS_CH = 8'h20;
    parameter [11:0] TL_CREDITS_NPD = 12'h028;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h198;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
    parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_MODE_ENABLE = "FALSE";
    parameter TL_PF_ENABLE_REG = "FALSE";
    parameter TL_TAG_MGMT_ENABLE = "TRUE";
    parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
    parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF0_PM_CAP_ID = 8'h01;
    parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
    parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF0_TPHR_CAP_ENABLE = "FALSE";
    parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF1_PM_CAP_ID = 8'h01;
    parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
    parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF1_TPHR_CAP_ENABLE = "FALSE";
    parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF2_PM_CAP_ID = 8'h01;
    parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
    parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF2_TPHR_CAP_ENABLE = "FALSE";
    parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF3_PM_CAP_ID = 8'h01;
    parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
    parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF3_TPHR_CAP_ENABLE = "FALSE";
    parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF4_PM_CAP_ID = 8'h01;
    parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
    parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF4_TPHR_CAP_ENABLE = "FALSE";
    parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF5_PM_CAP_ID = 8'h01;
    parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
    parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF5_TPHR_CAP_ENABLE = "FALSE";
    parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output CFGEXTREADRECEIVED;
    output CFGEXTWRITERECEIVED;
    output CFGHOTRESETOUT;
    output CFGINPUTUPDATEDONE;
    output CFGINTERRUPTAOUTPUT;
    output CFGINTERRUPTBOUTPUT;
    output CFGINTERRUPTCOUTPUT;
    output CFGINTERRUPTDOUTPUT;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output CFGINTERRUPTMSISENT;
    output CFGINTERRUPTMSIXFAIL;
    output CFGINTERRUPTMSIXSENT;
    output CFGINTERRUPTSENT;
    output CFGLOCALERROR;
    output CFGLTRENABLE;
    output CFGMCUPDATEDONE;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output CFGMSGTRANSMITDONE;
    output CFGPERFUNCTIONUPDATEDONE;
    output CFGPHYLINKDOWN;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output CFGTPHSTTREADENABLE;
    output CFGTPHSTTWRITEENABLE;
    output DRPRDY;
    output MAXISCQTLAST;
    output MAXISCQTVALID;
    output MAXISRCTLAST;
    output MAXISRCTVALID;
    output PCIERQSEQNUMVLD;
    output PCIERQTAGVLD;
    output PIPERX0POLARITY;
    output PIPERX1POLARITY;
    output PIPERX2POLARITY;
    output PIPERX3POLARITY;
    output PIPERX4POLARITY;
    output PIPERX5POLARITY;
    output PIPERX6POLARITY;
    output PIPERX7POLARITY;
    output PIPETX0COMPLIANCE;
    output PIPETX0DATAVALID;
    output PIPETX0ELECIDLE;
    output PIPETX0STARTBLOCK;
    output PIPETX1COMPLIANCE;
    output PIPETX1DATAVALID;
    output PIPETX1ELECIDLE;
    output PIPETX1STARTBLOCK;
    output PIPETX2COMPLIANCE;
    output PIPETX2DATAVALID;
    output PIPETX2ELECIDLE;
    output PIPETX2STARTBLOCK;
    output PIPETX3COMPLIANCE;
    output PIPETX3DATAVALID;
    output PIPETX3ELECIDLE;
    output PIPETX3STARTBLOCK;
    output PIPETX4COMPLIANCE;
    output PIPETX4DATAVALID;
    output PIPETX4ELECIDLE;
    output PIPETX4STARTBLOCK;
    output PIPETX5COMPLIANCE;
    output PIPETX5DATAVALID;
    output PIPETX5ELECIDLE;
    output PIPETX5STARTBLOCK;
    output PIPETX6COMPLIANCE;
    output PIPETX6DATAVALID;
    output PIPETX6ELECIDLE;
    output PIPETX6STARTBLOCK;
    output PIPETX7COMPLIANCE;
    output PIPETX7DATAVALID;
    output PIPETX7ELECIDLE;
    output PIPETX7STARTBLOCK;
    output PIPETXDEEMPH;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [11:0] CFGFCCPLD;
    output [11:0] CFGFCNPD;
    output [11:0] CFGFCPD;
    output [11:0] CFGVFSTATUS;
    output [143:0] MIREPLAYRAMWRITEDATA;
    output [143:0] MIREQUESTRAMWRITEDATA;
    output [15:0] CFGPERFUNCSTATUSDATA;
    output [15:0] DBGDATAOUT;
    output [15:0] DRPDO;
    output [17:0] CFGVFPOWERSTATE;
    output [17:0] CFGVFTPHSTMODE;
    output [1:0] CFGDPASUBSTATECHANGE;
    output [1:0] CFGFLRINPROCESS;
    output [1:0] CFGINTERRUPTMSIENABLE;
    output [1:0] CFGINTERRUPTMSIXENABLE;
    output [1:0] CFGINTERRUPTMSIXMASK;
    output [1:0] CFGLINKPOWERSTATE;
    output [1:0] CFGOBFFENABLE;
    output [1:0] CFGPHYLINKSTATUS;
    output [1:0] CFGRCBSTATUS;
    output [1:0] CFGTPHREQUESTERENABLE;
    output [1:0] MIREPLAYRAMREADENABLE;
    output [1:0] MIREPLAYRAMWRITEENABLE;
    output [1:0] PCIERQTAGAV;
    output [1:0] PCIETFCNPDAV;
    output [1:0] PCIETFCNPHAV;
    output [1:0] PIPERX0EQCONTROL;
    output [1:0] PIPERX1EQCONTROL;
    output [1:0] PIPERX2EQCONTROL;
    output [1:0] PIPERX3EQCONTROL;
    output [1:0] PIPERX4EQCONTROL;
    output [1:0] PIPERX5EQCONTROL;
    output [1:0] PIPERX6EQCONTROL;
    output [1:0] PIPERX7EQCONTROL;
    output [1:0] PIPETX0CHARISK;
    output [1:0] PIPETX0EQCONTROL;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX0SYNCHEADER;
    output [1:0] PIPETX1CHARISK;
    output [1:0] PIPETX1EQCONTROL;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX1SYNCHEADER;
    output [1:0] PIPETX2CHARISK;
    output [1:0] PIPETX2EQCONTROL;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX2SYNCHEADER;
    output [1:0] PIPETX3CHARISK;
    output [1:0] PIPETX3EQCONTROL;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX3SYNCHEADER;
    output [1:0] PIPETX4CHARISK;
    output [1:0] PIPETX4EQCONTROL;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX4SYNCHEADER;
    output [1:0] PIPETX5CHARISK;
    output [1:0] PIPETX5EQCONTROL;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX5SYNCHEADER;
    output [1:0] PIPETX6CHARISK;
    output [1:0] PIPETX6EQCONTROL;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX6SYNCHEADER;
    output [1:0] PIPETX7CHARISK;
    output [1:0] PIPETX7EQCONTROL;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PIPETX7SYNCHEADER;
    output [1:0] PIPETXRATE;
    output [1:0] PLEQPHASE;
    output [255:0] MAXISCQTDATA;
    output [255:0] MAXISRCTDATA;
    output [2:0] CFGCURRENTSPEED;
    output [2:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [2:0] CFGTPHFUNCTIONNUM;
    output [2:0] PIPERX0EQPRESET;
    output [2:0] PIPERX1EQPRESET;
    output [2:0] PIPERX2EQPRESET;
    output [2:0] PIPERX3EQPRESET;
    output [2:0] PIPERX4EQPRESET;
    output [2:0] PIPERX5EQPRESET;
    output [2:0] PIPERX6EQPRESET;
    output [2:0] PIPERX7EQPRESET;
    output [2:0] PIPETXMARGIN;
    output [31:0] CFGEXTWRITEDATA;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [31:0] CFGMGMTREADDATA;
    output [31:0] CFGTPHSTTWRITEDATA;
    output [31:0] PIPETX0DATA;
    output [31:0] PIPETX1DATA;
    output [31:0] PIPETX2DATA;
    output [31:0] PIPETX3DATA;
    output [31:0] PIPETX4DATA;
    output [31:0] PIPETX5DATA;
    output [31:0] PIPETX6DATA;
    output [31:0] PIPETX7DATA;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [3:0] CFGNEGOTIATEDWIDTH;
    output [3:0] CFGTPHSTTWRITEBYTEVALID;
    output [3:0] MICOMPLETIONRAMREADENABLEL;
    output [3:0] MICOMPLETIONRAMREADENABLEU;
    output [3:0] MICOMPLETIONRAMWRITEENABLEL;
    output [3:0] MICOMPLETIONRAMWRITEENABLEU;
    output [3:0] MIREQUESTRAMREADENABLE;
    output [3:0] MIREQUESTRAMWRITEENABLE;
    output [3:0] PCIERQSEQNUM;
    output [3:0] PIPERX0EQLPTXPRESET;
    output [3:0] PIPERX1EQLPTXPRESET;
    output [3:0] PIPERX2EQLPTXPRESET;
    output [3:0] PIPERX3EQLPTXPRESET;
    output [3:0] PIPERX4EQLPTXPRESET;
    output [3:0] PIPERX5EQLPTXPRESET;
    output [3:0] PIPERX6EQLPTXPRESET;
    output [3:0] PIPERX7EQLPTXPRESET;
    output [3:0] PIPETX0EQPRESET;
    output [3:0] PIPETX1EQPRESET;
    output [3:0] PIPETX2EQPRESET;
    output [3:0] PIPETX3EQPRESET;
    output [3:0] PIPETX4EQPRESET;
    output [3:0] PIPETX5EQPRESET;
    output [3:0] PIPETX6EQPRESET;
    output [3:0] PIPETX7EQPRESET;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output [4:0] CFGTPHSTTADDRESS;
    output [5:0] CFGFUNCTIONPOWERSTATE;
    output [5:0] CFGINTERRUPTMSIMMENABLE;
    output [5:0] CFGINTERRUPTMSIVFENABLE;
    output [5:0] CFGINTERRUPTMSIXVFENABLE;
    output [5:0] CFGINTERRUPTMSIXVFMASK;
    output [5:0] CFGLTSSMSTATE;
    output [5:0] CFGTPHSTMODE;
    output [5:0] CFGVFFLRINPROCESS;
    output [5:0] CFGVFTPHREQUESTERENABLE;
    output [5:0] PCIECQNPREQCOUNT;
    output [5:0] PCIERQTAG;
    output [5:0] PIPERX0EQLPLFFS;
    output [5:0] PIPERX1EQLPLFFS;
    output [5:0] PIPERX2EQLPLFFS;
    output [5:0] PIPERX3EQLPLFFS;
    output [5:0] PIPERX4EQLPLFFS;
    output [5:0] PIPERX5EQLPLFFS;
    output [5:0] PIPERX6EQLPLFFS;
    output [5:0] PIPERX7EQLPLFFS;
    output [5:0] PIPETX0EQDEEMPH;
    output [5:0] PIPETX1EQDEEMPH;
    output [5:0] PIPETX2EQDEEMPH;
    output [5:0] PIPETX3EQDEEMPH;
    output [5:0] PIPETX4EQDEEMPH;
    output [5:0] PIPETX5EQDEEMPH;
    output [5:0] PIPETX6EQDEEMPH;
    output [5:0] PIPETX7EQDEEMPH;
    output [71:0] MICOMPLETIONRAMWRITEDATAL;
    output [71:0] MICOMPLETIONRAMWRITEDATAU;
    output [74:0] MAXISRCTUSER;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output [7:0] CFGFCCPLH;
    output [7:0] CFGFCNPH;
    output [7:0] CFGFCPH;
    output [7:0] CFGFUNCTIONSTATUS;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [7:0] MAXISCQTKEEP;
    output [7:0] MAXISRCTKEEP;
    output [7:0] PLGEN3PCSRXSLIDE;
    output [84:0] MAXISCQTUSER;
    output [8:0] MIREPLAYRAMADDRESS;
    output [8:0] MIREQUESTRAMREADADDRESSA;
    output [8:0] MIREQUESTRAMREADADDRESSB;
    output [8:0] MIREQUESTRAMWRITEADDRESSA;
    output [8:0] MIREQUESTRAMWRITEADDRESSB;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [9:0] MICOMPLETIONRAMREADADDRESSAL;
    output [9:0] MICOMPLETIONRAMREADADDRESSAU;
    output [9:0] MICOMPLETIONRAMREADADDRESSBL;
    output [9:0] MICOMPLETIONRAMREADADDRESSBU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;
    input CFGCONFIGSPACEENABLE;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input CFGEXTREADDATAVALID;
    input CFGHOTRESETIN;
    input CFGINPUTUPDATEREQUEST;
    input CFGINTERRUPTMSITPHPRESENT;
    input CFGINTERRUPTMSIXINT;
    input CFGLINKTRAININGENABLE;
    input CFGMCUPDATEREQUEST;
    input CFGMGMTREAD;
    input CFGMGMTTYPE1CFGREGACCESS;
    input CFGMGMTWRITE;
    input CFGMSGTRANSMIT;
    input CFGPERFUNCTIONOUTPUTREQUEST;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input CFGTPHSTTREADDATAVALID;
    input CORECLK;
    input CORECLKMICOMPLETIONRAML;
    input CORECLKMICOMPLETIONRAMU;
    input CORECLKMIREPLAYRAM;
    input CORECLKMIREQUESTRAM;
    input DRPCLK;
    input DRPEN;
    input DRPWE;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input PCIECQNPREQ;
    input PIPECLK;
    input PIPERESETN;
    input PIPERX0DATAVALID;
    input PIPERX0ELECIDLE;
    input PIPERX0EQDONE;
    input PIPERX0EQLPADAPTDONE;
    input PIPERX0EQLPLFFSSEL;
    input PIPERX0PHYSTATUS;
    input PIPERX0STARTBLOCK;
    input PIPERX0VALID;
    input PIPERX1DATAVALID;
    input PIPERX1ELECIDLE;
    input PIPERX1EQDONE;
    input PIPERX1EQLPADAPTDONE;
    input PIPERX1EQLPLFFSSEL;
    input PIPERX1PHYSTATUS;
    input PIPERX1STARTBLOCK;
    input PIPERX1VALID;
    input PIPERX2DATAVALID;
    input PIPERX2ELECIDLE;
    input PIPERX2EQDONE;
    input PIPERX2EQLPADAPTDONE;
    input PIPERX2EQLPLFFSSEL;
    input PIPERX2PHYSTATUS;
    input PIPERX2STARTBLOCK;
    input PIPERX2VALID;
    input PIPERX3DATAVALID;
    input PIPERX3ELECIDLE;
    input PIPERX3EQDONE;
    input PIPERX3EQLPADAPTDONE;
    input PIPERX3EQLPLFFSSEL;
    input PIPERX3PHYSTATUS;
    input PIPERX3STARTBLOCK;
    input PIPERX3VALID;
    input PIPERX4DATAVALID;
    input PIPERX4ELECIDLE;
    input PIPERX4EQDONE;
    input PIPERX4EQLPADAPTDONE;
    input PIPERX4EQLPLFFSSEL;
    input PIPERX4PHYSTATUS;
    input PIPERX4STARTBLOCK;
    input PIPERX4VALID;
    input PIPERX5DATAVALID;
    input PIPERX5ELECIDLE;
    input PIPERX5EQDONE;
    input PIPERX5EQLPADAPTDONE;
    input PIPERX5EQLPLFFSSEL;
    input PIPERX5PHYSTATUS;
    input PIPERX5STARTBLOCK;
    input PIPERX5VALID;
    input PIPERX6DATAVALID;
    input PIPERX6ELECIDLE;
    input PIPERX6EQDONE;
    input PIPERX6EQLPADAPTDONE;
    input PIPERX6EQLPLFFSSEL;
    input PIPERX6PHYSTATUS;
    input PIPERX6STARTBLOCK;
    input PIPERX6VALID;
    input PIPERX7DATAVALID;
    input PIPERX7ELECIDLE;
    input PIPERX7EQDONE;
    input PIPERX7EQLPADAPTDONE;
    input PIPERX7EQLPLFFSSEL;
    input PIPERX7PHYSTATUS;
    input PIPERX7STARTBLOCK;
    input PIPERX7VALID;
    input PIPETX0EQDONE;
    input PIPETX1EQDONE;
    input PIPETX2EQDONE;
    input PIPETX3EQDONE;
    input PIPETX4EQDONE;
    input PIPETX5EQDONE;
    input PIPETX6EQDONE;
    input PIPETX7EQDONE;
    input PLDISABLESCRAMBLER;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN3PCSDISABLE;
    input RECCLK;
    input RESETN;
    input SAXISCCTLAST;
    input SAXISCCTVALID;
    input SAXISRQTLAST;
    input SAXISRQTVALID;
    input USERCLK;
    input [10:0] DRPADDR;
    input [143:0] MICOMPLETIONRAMREADDATA;
    input [143:0] MIREPLAYRAMREADDATA;
    input [143:0] MIREQUESTRAMREADDATA;
    input [15:0] CFGDEVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [15:0] CFGVENDID;
    input [15:0] DRPDI;
    input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
    input [17:0] PIPETX0EQCOEFF;
    input [17:0] PIPETX1EQCOEFF;
    input [17:0] PIPETX2EQCOEFF;
    input [17:0] PIPETX3EQCOEFF;
    input [17:0] PIPETX4EQCOEFF;
    input [17:0] PIPETX5EQCOEFF;
    input [17:0] PIPETX6EQCOEFF;
    input [17:0] PIPETX7EQCOEFF;
    input [18:0] CFGMGMTADDR;
    input [1:0] CFGFLRDONE;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [1:0] CFGINTERRUPTPENDING;
    input [1:0] PIPERX0CHARISK;
    input [1:0] PIPERX0SYNCHEADER;
    input [1:0] PIPERX1CHARISK;
    input [1:0] PIPERX1SYNCHEADER;
    input [1:0] PIPERX2CHARISK;
    input [1:0] PIPERX2SYNCHEADER;
    input [1:0] PIPERX3CHARISK;
    input [1:0] PIPERX3SYNCHEADER;
    input [1:0] PIPERX4CHARISK;
    input [1:0] PIPERX4SYNCHEADER;
    input [1:0] PIPERX5CHARISK;
    input [1:0] PIPERX5SYNCHEADER;
    input [1:0] PIPERX6CHARISK;
    input [1:0] PIPERX6SYNCHEADER;
    input [1:0] PIPERX7CHARISK;
    input [1:0] PIPERX7SYNCHEADER;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input [255:0] SAXISCCTDATA;
    input [255:0] SAXISRQTDATA;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [2:0] CFGFCSEL;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [2:0] CFGPERFUNCSTATUSCONTROL;
    input [2:0] CFGPERFUNCTIONNUMBER;
    input [2:0] PIPERX0STATUS;
    input [2:0] PIPERX1STATUS;
    input [2:0] PIPERX2STATUS;
    input [2:0] PIPERX3STATUS;
    input [2:0] PIPERX4STATUS;
    input [2:0] PIPERX5STATUS;
    input [2:0] PIPERX6STATUS;
    input [2:0] PIPERX7STATUS;
    input [31:0] CFGEXTREADDATA;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input [31:0] CFGMGMTWRITEDATA;
    input [31:0] CFGMSGTRANSMITDATA;
    input [31:0] CFGTPHSTTREADDATA;
    input [31:0] PIPERX0DATA;
    input [31:0] PIPERX1DATA;
    input [31:0] PIPERX2DATA;
    input [31:0] PIPERX3DATA;
    input [31:0] PIPERX4DATA;
    input [31:0] PIPERX5DATA;
    input [31:0] PIPERX6DATA;
    input [31:0] PIPERX7DATA;
    input [32:0] SAXISCCTUSER;
    input [3:0] CFGINTERRUPTINT;
    input [3:0] CFGINTERRUPTMSISELECT;
    input [3:0] CFGMGMTBYTEENABLE;
    input [4:0] CFGDSDEVICENUMBER;
    input [59:0] SAXISRQTUSER;
    input [5:0] CFGVFFLRDONE;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input [63:0] CFGDSN;
    input [63:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [7:0] CFGDSBUSNUMBER;
    input [7:0] CFGDSPORTNUMBER;
    input [7:0] CFGREVID;
    input [7:0] PLGEN3PCSRXSYNCDONE;
    input [7:0] SAXISCCTKEEP;
    input [7:0] SAXISRQTKEEP;
    input [8:0] CFGINTERRUPTMSITPHSTTAG;
endmodule

module PCIE_3_1 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
    parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
    parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE = "FALSE";
    parameter DEBUG_PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
    parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF0_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_BIST_REGISTER = 8'h00;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter [15:0] PF0_DEVICE_ID = 16'h0000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF0_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
    parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF0_PB_CAP_VER = 4'h1;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter PF0_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF0_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF0_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF0_RBAR_NUM = 3'h1;
    parameter [7:0] PF0_REVISION_ID = 8'h00;
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF1_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_BIST_REGISTER = 8'h00;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [15:0] PF1_DEVICE_ID = 16'h0000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF1_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
    parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF1_PB_CAP_VER = 4'h1;
    parameter [7:0] PF1_PM_CAP_ID = 8'h01;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
    parameter PF1_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF1_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF1_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF1_RBAR_NUM = 3'h1;
    parameter [7:0] PF1_REVISION_ID = 8'h00;
    parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
    parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF1_TPHR_CAP_ENABLE = "FALSE";
    parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
    parameter PF2_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF2_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF2_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_BIST_REGISTER = 8'h00;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [15:0] PF2_DEVICE_ID = 16'h0000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF2_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF2_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF2_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF2_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF2_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF2_PB_CAP_NEXTPTR = 12'h000;
    parameter PF2_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF2_PB_CAP_VER = 4'h1;
    parameter [7:0] PF2_PM_CAP_ID = 8'h01;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF2_PM_CAP_VER_ID = 3'h3;
    parameter PF2_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF2_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF2_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF2_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF2_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF2_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF2_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF2_RBAR_NUM = 3'h1;
    parameter [7:0] PF2_REVISION_ID = 8'h00;
    parameter [4:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF2_SUBSYSTEM_ID = 16'h0000;
    parameter PF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF2_TPHR_CAP_ENABLE = "FALSE";
    parameter PF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF2_TPHR_CAP_VER = 4'h1;
    parameter PF3_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
    parameter PF3_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [5:0] PF3_BAR1_APERTURE_SIZE = 6'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_BIST_REGISTER = 8'h00;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h50;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [15:0] PF3_DEVICE_ID = 16'h0000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DPA_CAP_NEXTPTR = 12'h000;
    parameter [4:0] PF3_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
    parameter PF3_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
    parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
    parameter [3:0] PF3_DPA_CAP_VER = 4'h1;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [7:0] PF3_INTERRUPT_LINE = 8'h00;
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D1 = 32'h00000000;
    parameter [31:0] PF3_PB_CAP_DATA_REG_D3HOT = 32'h00000000;
    parameter [11:0] PF3_PB_CAP_NEXTPTR = 12'h000;
    parameter PF3_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
    parameter [3:0] PF3_PB_CAP_VER = 4'h1;
    parameter [7:0] PF3_PM_CAP_ID = 8'h01;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] PF3_PM_CAP_VER_ID = 3'h3;
    parameter PF3_RBAR_CAP_ENABLE = "FALSE";
    parameter [11:0] PF3_RBAR_CAP_NEXTPTR = 12'h000;
    parameter [19:0] PF3_RBAR_CAP_SIZE0 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE1 = 20'h00000;
    parameter [19:0] PF3_RBAR_CAP_SIZE2 = 20'h00000;
    parameter [3:0] PF3_RBAR_CAP_VER = 4'h1;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX0 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX1 = 3'h0;
    parameter [2:0] PF3_RBAR_CONTROL_INDEX2 = 3'h0;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE0 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE1 = 5'h00;
    parameter [4:0] PF3_RBAR_CONTROL_SIZE2 = 5'h00;
    parameter [2:0] PF3_RBAR_NUM = 3'h1;
    parameter [7:0] PF3_REVISION_ID = 8'h00;
    parameter [4:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [4:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [15:0] PF3_SUBSYSTEM_ID = 16'h0000;
    parameter PF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF3_TPHR_CAP_ENABLE = "FALSE";
    parameter PF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF3_TPHR_CAP_VER = 4'h1;
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP = "TRUE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_SCRAMBLING = "FALSE";
    parameter PL_DISABLE_SYNC_HEADER_FRAMING_ERROR = "FALSE";
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
    parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
    parameter [2:0] PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT = 3'h3;
    parameter [3:0] PL_EQ_DEFAULT_GEN3_TX_PRESET = 4'h4;
    parameter PL_EQ_PHASE01_RX_ADAPT = "FALSE";
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
    parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
    parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
    parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
    parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
    parameter integer PL_N_FTS_GEN1 = 255;
    parameter integer PL_N_FTS_GEN2 = 255;
    parameter integer PL_N_FTS_GEN3 = 255;
    parameter PL_REPORT_ALL_PHY_ERRORS = "TRUE";
    parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter integer SPARE_BIT0 = 0;
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter integer SPARE_BIT3 = 0;
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter SRIOV_CAP_ENABLE = "FALSE";
    parameter TL_COMPLETION_RAM_SIZE_16K = "TRUE";
    parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [11:0] TL_CREDITS_CD = 12'h3E0;
    parameter [7:0] TL_CREDITS_CH = 8'h20;
    parameter [11:0] TL_CREDITS_NPD = 12'h028;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h198;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
    parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter TL_LEGACY_MODE_ENABLE = "FALSE";
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TWO_LAYER_MODE_DLCMSM_ENABLE = "TRUE";
    parameter TWO_LAYER_MODE_ENABLE = "FALSE";
    parameter TWO_LAYER_MODE_WIDTH_256 = "TRUE";
    parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
    parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF0_PM_CAP_ID = 8'h01;
    parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
    parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF0_TPHR_CAP_ENABLE = "FALSE";
    parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF1_PM_CAP_ID = 8'h01;
    parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
    parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF1_TPHR_CAP_ENABLE = "FALSE";
    parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF2_PM_CAP_ID = 8'h01;
    parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
    parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF2_TPHR_CAP_ENABLE = "FALSE";
    parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF3_PM_CAP_ID = 8'h01;
    parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
    parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF3_TPHR_CAP_ENABLE = "FALSE";
    parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF4_PM_CAP_ID = 8'h01;
    parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
    parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF4_TPHR_CAP_ENABLE = "FALSE";
    parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF5_PM_CAP_ID = 8'h01;
    parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
    parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF5_TPHR_CAP_ENABLE = "FALSE";
    parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF6_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF6_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF6_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF6_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF6_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF6_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF6_PM_CAP_ID = 8'h01;
    parameter [7:0] VF6_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF6_PM_CAP_VER_ID = 3'h3;
    parameter VF6_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF6_TPHR_CAP_ENABLE = "FALSE";
    parameter VF6_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF6_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF6_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF6_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF6_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF6_TPHR_CAP_VER = 4'h1;
    parameter [11:0] VF7_ARI_CAP_NEXTPTR = 12'h000;
    parameter integer VF7_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VF7_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VF7_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VF7_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer VF7_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] VF7_PM_CAP_ID = 8'h01;
    parameter [7:0] VF7_PM_CAP_NEXTPTR = 8'h00;
    parameter [2:0] VF7_PM_CAP_VER_ID = 3'h3;
    parameter VF7_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter VF7_TPHR_CAP_ENABLE = "FALSE";
    parameter VF7_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] VF7_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VF7_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] VF7_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] VF7_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] VF7_TPHR_CAP_VER = 4'h1;
    output [2:0] CFGCURRENTSPEED;
    output [3:0] CFGDPASUBSTATECHANGE;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [7:0] CFGINTERRUPTMSIVFENABLE;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output CFGINTERRUPTMSIXFAIL;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXSENT;
    output [7:0] CFGINTERRUPTMSIXVFENABLE;
    output [7:0] CFGINTERRUPTMSIXVFMASK;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output CFGLOCALERROR;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [2:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [3:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output [15:0] CFGPERFUNCSTATUSDATA;
    output CFGPERFUNCTIONUPDATEDONE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [3:0] CFGTPHFUNCTIONNUM;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [4:0] CFGTPHSTTADDRESS;
    output CFGTPHSTTREADENABLE;
    output [3:0] CFGTPHSTTWRITEBYTEVALID;
    output [31:0] CFGTPHSTTWRITEDATA;
    output CFGTPHSTTWRITEENABLE;
    output [7:0] CFGVFFLRINPROCESS;
    output [23:0] CFGVFPOWERSTATE;
    output [15:0] CFGVFSTATUS;
    output [7:0] CFGVFTPHREQUESTERENABLE;
    output [23:0] CFGVFTPHSTMODE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [15:0] DBGDATAOUT;
    output DBGMCAPCSB;
    output [31:0] DBGMCAPDATA;
    output DBGMCAPEOS;
    output DBGMCAPERROR;
    output DBGMCAPMODE;
    output DBGMCAPRDATAVALID;
    output DBGMCAPRDWRB;
    output DBGMCAPRESET;
    output DBGPLDATABLOCKRECEIVEDAFTEREDS;
    output DBGPLGEN3FRAMINGERRORDETECTED;
    output DBGPLGEN3SYNCHEADERERRORDETECTED;
    output [7:0] DBGPLINFERREDRXELECTRICALIDLE;
    output [15:0] DRPDO;
    output DRPRDY;
    output LL2LMMASTERTLPSENT0;
    output LL2LMMASTERTLPSENT1;
    output [3:0] LL2LMMASTERTLPSENTTLPID0;
    output [3:0] LL2LMMASTERTLPSENTTLPID1;
    output [255:0] LL2LMMAXISRXTDATA;
    output [17:0] LL2LMMAXISRXTUSER;
    output [7:0] LL2LMMAXISRXTVALID;
    output [7:0] LL2LMSAXISTXTREADY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [84:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [9:0] MICOMPLETIONRAMREADADDRESSAL;
    output [9:0] MICOMPLETIONRAMREADADDRESSAU;
    output [9:0] MICOMPLETIONRAMREADADDRESSBL;
    output [9:0] MICOMPLETIONRAMREADADDRESSBU;
    output [3:0] MICOMPLETIONRAMREADENABLEL;
    output [3:0] MICOMPLETIONRAMREADENABLEU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
    output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;
    output [71:0] MICOMPLETIONRAMWRITEDATAL;
    output [71:0] MICOMPLETIONRAMWRITEDATAU;
    output [3:0] MICOMPLETIONRAMWRITEENABLEL;
    output [3:0] MICOMPLETIONRAMWRITEENABLEU;
    output [8:0] MIREPLAYRAMADDRESS;
    output [1:0] MIREPLAYRAMREADENABLE;
    output [143:0] MIREPLAYRAMWRITEDATA;
    output [1:0] MIREPLAYRAMWRITEENABLE;
    output [8:0] MIREQUESTRAMREADADDRESSA;
    output [8:0] MIREQUESTRAMREADADDRESSB;
    output [3:0] MIREQUESTRAMREADENABLE;
    output [8:0] MIREQUESTRAMWRITEADDRESSA;
    output [8:0] MIREQUESTRAMWRITEADDRESSB;
    output [143:0] MIREQUESTRAMWRITEDATA;
    output [3:0] MIREQUESTRAMWRITEENABLE;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [3:0] PCIERQSEQNUM;
    output PCIERQSEQNUMVLD;
    output [5:0] PCIERQTAG;
    output [1:0] PCIERQTAGAV;
    output PCIERQTAGVLD;
    output [1:0] PCIETFCNPDAV;
    output [1:0] PCIETFCNPHAV;
    output [1:0] PIPERX0EQCONTROL;
    output [5:0] PIPERX0EQLPLFFS;
    output [3:0] PIPERX0EQLPTXPRESET;
    output [2:0] PIPERX0EQPRESET;
    output PIPERX0POLARITY;
    output [1:0] PIPERX1EQCONTROL;
    output [5:0] PIPERX1EQLPLFFS;
    output [3:0] PIPERX1EQLPTXPRESET;
    output [2:0] PIPERX1EQPRESET;
    output PIPERX1POLARITY;
    output [1:0] PIPERX2EQCONTROL;
    output [5:0] PIPERX2EQLPLFFS;
    output [3:0] PIPERX2EQLPTXPRESET;
    output [2:0] PIPERX2EQPRESET;
    output PIPERX2POLARITY;
    output [1:0] PIPERX3EQCONTROL;
    output [5:0] PIPERX3EQLPLFFS;
    output [3:0] PIPERX3EQLPTXPRESET;
    output [2:0] PIPERX3EQPRESET;
    output PIPERX3POLARITY;
    output [1:0] PIPERX4EQCONTROL;
    output [5:0] PIPERX4EQLPLFFS;
    output [3:0] PIPERX4EQLPTXPRESET;
    output [2:0] PIPERX4EQPRESET;
    output PIPERX4POLARITY;
    output [1:0] PIPERX5EQCONTROL;
    output [5:0] PIPERX5EQLPLFFS;
    output [3:0] PIPERX5EQLPTXPRESET;
    output [2:0] PIPERX5EQPRESET;
    output PIPERX5POLARITY;
    output [1:0] PIPERX6EQCONTROL;
    output [5:0] PIPERX6EQLPLFFS;
    output [3:0] PIPERX6EQLPTXPRESET;
    output [2:0] PIPERX6EQPRESET;
    output PIPERX6POLARITY;
    output [1:0] PIPERX7EQCONTROL;
    output [5:0] PIPERX7EQLPLFFS;
    output [3:0] PIPERX7EQLPTXPRESET;
    output [2:0] PIPERX7EQPRESET;
    output PIPERX7POLARITY;
    output [1:0] PIPETX0CHARISK;
    output PIPETX0COMPLIANCE;
    output [31:0] PIPETX0DATA;
    output PIPETX0DATAVALID;
    output PIPETX0DEEMPH;
    output PIPETX0ELECIDLE;
    output [1:0] PIPETX0EQCONTROL;
    output [5:0] PIPETX0EQDEEMPH;
    output [3:0] PIPETX0EQPRESET;
    output [2:0] PIPETX0MARGIN;
    output [1:0] PIPETX0POWERDOWN;
    output [1:0] PIPETX0RATE;
    output PIPETX0RCVRDET;
    output PIPETX0RESET;
    output PIPETX0STARTBLOCK;
    output PIPETX0SWING;
    output [1:0] PIPETX0SYNCHEADER;
    output [1:0] PIPETX1CHARISK;
    output PIPETX1COMPLIANCE;
    output [31:0] PIPETX1DATA;
    output PIPETX1DATAVALID;
    output PIPETX1DEEMPH;
    output PIPETX1ELECIDLE;
    output [1:0] PIPETX1EQCONTROL;
    output [5:0] PIPETX1EQDEEMPH;
    output [3:0] PIPETX1EQPRESET;
    output [2:0] PIPETX1MARGIN;
    output [1:0] PIPETX1POWERDOWN;
    output [1:0] PIPETX1RATE;
    output PIPETX1RCVRDET;
    output PIPETX1RESET;
    output PIPETX1STARTBLOCK;
    output PIPETX1SWING;
    output [1:0] PIPETX1SYNCHEADER;
    output [1:0] PIPETX2CHARISK;
    output PIPETX2COMPLIANCE;
    output [31:0] PIPETX2DATA;
    output PIPETX2DATAVALID;
    output PIPETX2DEEMPH;
    output PIPETX2ELECIDLE;
    output [1:0] PIPETX2EQCONTROL;
    output [5:0] PIPETX2EQDEEMPH;
    output [3:0] PIPETX2EQPRESET;
    output [2:0] PIPETX2MARGIN;
    output [1:0] PIPETX2POWERDOWN;
    output [1:0] PIPETX2RATE;
    output PIPETX2RCVRDET;
    output PIPETX2RESET;
    output PIPETX2STARTBLOCK;
    output PIPETX2SWING;
    output [1:0] PIPETX2SYNCHEADER;
    output [1:0] PIPETX3CHARISK;
    output PIPETX3COMPLIANCE;
    output [31:0] PIPETX3DATA;
    output PIPETX3DATAVALID;
    output PIPETX3DEEMPH;
    output PIPETX3ELECIDLE;
    output [1:0] PIPETX3EQCONTROL;
    output [5:0] PIPETX3EQDEEMPH;
    output [3:0] PIPETX3EQPRESET;
    output [2:0] PIPETX3MARGIN;
    output [1:0] PIPETX3POWERDOWN;
    output [1:0] PIPETX3RATE;
    output PIPETX3RCVRDET;
    output PIPETX3RESET;
    output PIPETX3STARTBLOCK;
    output PIPETX3SWING;
    output [1:0] PIPETX3SYNCHEADER;
    output [1:0] PIPETX4CHARISK;
    output PIPETX4COMPLIANCE;
    output [31:0] PIPETX4DATA;
    output PIPETX4DATAVALID;
    output PIPETX4DEEMPH;
    output PIPETX4ELECIDLE;
    output [1:0] PIPETX4EQCONTROL;
    output [5:0] PIPETX4EQDEEMPH;
    output [3:0] PIPETX4EQPRESET;
    output [2:0] PIPETX4MARGIN;
    output [1:0] PIPETX4POWERDOWN;
    output [1:0] PIPETX4RATE;
    output PIPETX4RCVRDET;
    output PIPETX4RESET;
    output PIPETX4STARTBLOCK;
    output PIPETX4SWING;
    output [1:0] PIPETX4SYNCHEADER;
    output [1:0] PIPETX5CHARISK;
    output PIPETX5COMPLIANCE;
    output [31:0] PIPETX5DATA;
    output PIPETX5DATAVALID;
    output PIPETX5DEEMPH;
    output PIPETX5ELECIDLE;
    output [1:0] PIPETX5EQCONTROL;
    output [5:0] PIPETX5EQDEEMPH;
    output [3:0] PIPETX5EQPRESET;
    output [2:0] PIPETX5MARGIN;
    output [1:0] PIPETX5POWERDOWN;
    output [1:0] PIPETX5RATE;
    output PIPETX5RCVRDET;
    output PIPETX5RESET;
    output PIPETX5STARTBLOCK;
    output PIPETX5SWING;
    output [1:0] PIPETX5SYNCHEADER;
    output [1:0] PIPETX6CHARISK;
    output PIPETX6COMPLIANCE;
    output [31:0] PIPETX6DATA;
    output PIPETX6DATAVALID;
    output PIPETX6DEEMPH;
    output PIPETX6ELECIDLE;
    output [1:0] PIPETX6EQCONTROL;
    output [5:0] PIPETX6EQDEEMPH;
    output [3:0] PIPETX6EQPRESET;
    output [2:0] PIPETX6MARGIN;
    output [1:0] PIPETX6POWERDOWN;
    output [1:0] PIPETX6RATE;
    output PIPETX6RCVRDET;
    output PIPETX6RESET;
    output PIPETX6STARTBLOCK;
    output PIPETX6SWING;
    output [1:0] PIPETX6SYNCHEADER;
    output [1:0] PIPETX7CHARISK;
    output PIPETX7COMPLIANCE;
    output [31:0] PIPETX7DATA;
    output PIPETX7DATAVALID;
    output PIPETX7DEEMPH;
    output PIPETX7ELECIDLE;
    output [1:0] PIPETX7EQCONTROL;
    output [5:0] PIPETX7EQDEEMPH;
    output [3:0] PIPETX7EQPRESET;
    output [2:0] PIPETX7MARGIN;
    output [1:0] PIPETX7POWERDOWN;
    output [1:0] PIPETX7RATE;
    output PIPETX7RCVRDET;
    output PIPETX7RESET;
    output PIPETX7STARTBLOCK;
    output PIPETX7SWING;
    output [1:0] PIPETX7SYNCHEADER;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] SPAREOUT;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVID;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [3:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [8:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [18:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTREAD;
    input CFGMGMTTYPE1CFGREGACCESS;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [2:0] CFGPERFUNCSTATUSCONTROL;
    input [3:0] CFGPERFUNCTIONNUMBER;
    input CFGPERFUNCTIONOUTPUTREQUEST;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVID;
    input [15:0] CFGSUBSYSID;
    input [15:0] CFGSUBSYSVENDID;
    input [31:0] CFGTPHSTTREADDATA;
    input CFGTPHSTTREADDATAVALID;
    input [15:0] CFGVENDID;
    input [7:0] CFGVFFLRDONE;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMICOMPLETIONRAML;
    input CORECLKMICOMPLETIONRAMU;
    input CORECLKMIREPLAYRAM;
    input CORECLKMIREQUESTRAM;
    input DBGCFGLOCALMGMTREGOVERRIDE;
    input [3:0] DBGDATASEL;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [13:0] LL2LMSAXISTXTUSER;
    input LL2LMSAXISTXTVALID;
    input [3:0] LL2LMTXTLPID0;
    input [3:0] LL2LMTXTLPID1;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [143:0] MICOMPLETIONRAMREADDATA;
    input [143:0] MIREPLAYRAMREADDATA;
    input [143:0] MIREQUESTRAMREADDATA;
    input PCIECQNPREQ;
    input PIPECLK;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX0CHARISK;
    input [31:0] PIPERX0DATA;
    input PIPERX0DATAVALID;
    input PIPERX0ELECIDLE;
    input PIPERX0EQDONE;
    input PIPERX0EQLPADAPTDONE;
    input PIPERX0EQLPLFFSSEL;
    input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
    input PIPERX0PHYSTATUS;
    input PIPERX0STARTBLOCK;
    input [2:0] PIPERX0STATUS;
    input [1:0] PIPERX0SYNCHEADER;
    input PIPERX0VALID;
    input [1:0] PIPERX1CHARISK;
    input [31:0] PIPERX1DATA;
    input PIPERX1DATAVALID;
    input PIPERX1ELECIDLE;
    input PIPERX1EQDONE;
    input PIPERX1EQLPADAPTDONE;
    input PIPERX1EQLPLFFSSEL;
    input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
    input PIPERX1PHYSTATUS;
    input PIPERX1STARTBLOCK;
    input [2:0] PIPERX1STATUS;
    input [1:0] PIPERX1SYNCHEADER;
    input PIPERX1VALID;
    input [1:0] PIPERX2CHARISK;
    input [31:0] PIPERX2DATA;
    input PIPERX2DATAVALID;
    input PIPERX2ELECIDLE;
    input PIPERX2EQDONE;
    input PIPERX2EQLPADAPTDONE;
    input PIPERX2EQLPLFFSSEL;
    input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
    input PIPERX2PHYSTATUS;
    input PIPERX2STARTBLOCK;
    input [2:0] PIPERX2STATUS;
    input [1:0] PIPERX2SYNCHEADER;
    input PIPERX2VALID;
    input [1:0] PIPERX3CHARISK;
    input [31:0] PIPERX3DATA;
    input PIPERX3DATAVALID;
    input PIPERX3ELECIDLE;
    input PIPERX3EQDONE;
    input PIPERX3EQLPADAPTDONE;
    input PIPERX3EQLPLFFSSEL;
    input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
    input PIPERX3PHYSTATUS;
    input PIPERX3STARTBLOCK;
    input [2:0] PIPERX3STATUS;
    input [1:0] PIPERX3SYNCHEADER;
    input PIPERX3VALID;
    input [1:0] PIPERX4CHARISK;
    input [31:0] PIPERX4DATA;
    input PIPERX4DATAVALID;
    input PIPERX4ELECIDLE;
    input PIPERX4EQDONE;
    input PIPERX4EQLPADAPTDONE;
    input PIPERX4EQLPLFFSSEL;
    input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
    input PIPERX4PHYSTATUS;
    input PIPERX4STARTBLOCK;
    input [2:0] PIPERX4STATUS;
    input [1:0] PIPERX4SYNCHEADER;
    input PIPERX4VALID;
    input [1:0] PIPERX5CHARISK;
    input [31:0] PIPERX5DATA;
    input PIPERX5DATAVALID;
    input PIPERX5ELECIDLE;
    input PIPERX5EQDONE;
    input PIPERX5EQLPADAPTDONE;
    input PIPERX5EQLPLFFSSEL;
    input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
    input PIPERX5PHYSTATUS;
    input PIPERX5STARTBLOCK;
    input [2:0] PIPERX5STATUS;
    input [1:0] PIPERX5SYNCHEADER;
    input PIPERX5VALID;
    input [1:0] PIPERX6CHARISK;
    input [31:0] PIPERX6DATA;
    input PIPERX6DATAVALID;
    input PIPERX6ELECIDLE;
    input PIPERX6EQDONE;
    input PIPERX6EQLPADAPTDONE;
    input PIPERX6EQLPLFFSSEL;
    input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
    input PIPERX6PHYSTATUS;
    input PIPERX6STARTBLOCK;
    input [2:0] PIPERX6STATUS;
    input [1:0] PIPERX6SYNCHEADER;
    input PIPERX6VALID;
    input [1:0] PIPERX7CHARISK;
    input [31:0] PIPERX7DATA;
    input PIPERX7DATAVALID;
    input PIPERX7ELECIDLE;
    input PIPERX7EQDONE;
    input PIPERX7EQLPADAPTDONE;
    input PIPERX7EQLPLFFSSEL;
    input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
    input PIPERX7PHYSTATUS;
    input PIPERX7STARTBLOCK;
    input [2:0] PIPERX7STATUS;
    input [1:0] PIPERX7SYNCHEADER;
    input PIPERX7VALID;
    input [17:0] PIPETX0EQCOEFF;
    input PIPETX0EQDONE;
    input [17:0] PIPETX1EQCOEFF;
    input PIPETX1EQDONE;
    input [17:0] PIPETX2EQCOEFF;
    input PIPETX2EQDONE;
    input [17:0] PIPETX3EQCOEFF;
    input PIPETX3EQDONE;
    input [17:0] PIPETX4EQCOEFF;
    input PIPETX4EQDONE;
    input [17:0] PIPETX5EQCOEFF;
    input PIPETX5EQDONE;
    input [17:0] PIPETX6EQCOEFF;
    input PIPETX6EQDONE;
    input [17:0] PIPETX7EQCOEFF;
    input PIPETX7EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [59:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input [31:0] SPAREIN;
    input USERCLK;
endmodule

module PCIE40E4 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AUTO_FLR_RESPONSE = "FALSE";
    parameter [1:0] AXISTEN_IF_CC_ALIGNMENT_MODE = 2'h0;
    parameter [23:0] AXISTEN_IF_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] AXISTEN_IF_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [1:0] AXISTEN_IF_CQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_CQ_EN_POISONED_MEM_WR = "FALSE";
    parameter AXISTEN_IF_ENABLE_256_TAGS = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE = "FALSE";
    parameter AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK = "TRUE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_EXT_512 = "FALSE";
    parameter AXISTEN_IF_EXT_512_CC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_CQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_LEGACY_MODE_ENABLE = "FALSE";
    parameter AXISTEN_IF_MSIX_FROM_RAM_PIPELINE = "FALSE";
    parameter AXISTEN_IF_MSIX_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_MSIX_TO_RAM_PIPELINE = "FALSE";
    parameter [1:0] AXISTEN_IF_RC_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter [1:0] AXISTEN_IF_RQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT = "FALSE";
    parameter AXISTEN_IF_TX_PARITY_EN = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CFG_BYPASS_MODE_ENABLE = "FALSE";
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [15:0] DEBUG_AXI4ST_SPARE = 16'h0000;
    parameter [7:0] DEBUG_AXIST_DISABLE_FEATURE_BIT = 8'h00;
    parameter [3:0] DEBUG_CAR_SPARE = 4'h0;
    parameter [15:0] DEBUG_CFG_SPARE = 16'h0000;
    parameter [15:0] DEBUG_LL_SPARE = 16'h0000;
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW = "FALSE";
    parameter DEBUG_PL_DISABLE_SCRAMBLING = "FALSE";
    parameter DEBUG_PL_SIM_RESET_LFSR = "FALSE";
    parameter [15:0] DEBUG_PL_SPARE = 16'h0000;
    parameter DEBUG_TL_DISABLE_FC_TIMEOUT = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [15:0] DEBUG_TL_SPARE = 16'h0000;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter DSN_CAP_ENABLE = "FALSE";
    parameter EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter HEADER_TYPE_OVERRIDE = "FALSE";
    parameter IS_SWITCH_PORT = "FALSE";
    parameter LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter LL_DISABLE_SCHED_TX_NAK = "FALSE";
    parameter LL_REPLAY_FROM_RAM_PIPELINE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter LL_REPLAY_TO_RAM_PIPELINE = "FALSE";
    parameter LL_RX_TLP_PARITY_GEN = "TRUE";
    parameter LL_TX_TLP_PARITY_CHK = "TRUE";
    parameter [15:0] LL_USER_SPARE = 16'h0000;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h250;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4 = 7;
    parameter [0:0] PF0_LINK_CONTROL_RCB = 1'h0;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [5:0] PF0_MSIX_VECTOR_COUNT = 6'h04;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter PL_CFG_STATE_ROBUSTNESS_ENABLE = "TRUE";
    parameter PL_DEEMPH_SOURCE_SELECT = "TRUE";
    parameter PL_DESKEW_ON_SKIP_IN_GEN12 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_LANE_REVERSAL = "FALSE";
    parameter [1:0] PL_DISABLE_LFSR_UPDATE_ON_SKP = 2'h0;
    parameter PL_DISABLE_RETRAIN_ON_EB_ERROR = "FALSE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter [15:0] PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR = 16'h0000;
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter [1:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK = 2'h0;
    parameter [1:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK = 2'h0;
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter [1:0] PL_EQ_BYPASS_PHASE23 = 2'h0;
    parameter [5:0] PL_EQ_DEFAULT_RX_PRESET_HINT = 6'h33;
    parameter [7:0] PL_EQ_DEFAULT_TX_PRESET = 8'h44;
    parameter PL_EQ_DISABLE_MISMATCH_CHECK = "TRUE";
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE0 = 2'h0;
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE1 = 2'h0;
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter PL_EQ_TX_8G_EQ_TS2_ENABLE = "FALSE";
    parameter PL_EXIT_LOOPBACK_ON_EI_ENTRY = "TRUE";
    parameter PL_INFER_EI_DISABLE_LPBK_ACTIVE = "TRUE";
    parameter PL_INFER_EI_DISABLE_REC_RC = "FALSE";
    parameter PL_INFER_EI_DISABLE_REC_SPD = "FALSE";
    parameter [31:0] PL_LANE0_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE10_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE11_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE12_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE13_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE14_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE15_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE1_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE2_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE3_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE4_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE5_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE6_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE7_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE8_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE9_EQ_CONTROL = 32'h00003F00;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_SPEED = 4'h4;
    parameter [4:0] PL_LINK_CAP_MAX_LINK_WIDTH = 5'h08;
    parameter integer PL_N_FTS = 255;
    parameter PL_QUIESCE_GUARANTEE_DISABLE = "FALSE";
    parameter PL_REDO_EQ_SOURCE_SELECT = "TRUE";
    parameter [7:0] PL_REPORT_ALL_PHY_ERRORS = 8'h00;
    parameter [1:0] PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN4 = 4'h0;
    parameter [1:0] PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN4 = 4'h0;
    parameter [1:0] PL_RX_L0S_EXIT_TO_RECOVERY = 2'h0;
    parameter [1:0] PL_SIM_FAST_LINK_TRAINING = 2'h0;
    parameter PL_SRIS_ENABLE = "FALSE";
    parameter [6:0] PL_SRIS_SKPOS_GEN_SPD_VEC = 7'h00;
    parameter [6:0] PL_SRIS_SKPOS_REC_SPD_VEC = 7'h00;
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PL_USER_SPARE = 16'h0000;
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h1500;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h003E8;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000100;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h00000;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0100;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter SPARE_BIT0 = "FALSE";
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter SPARE_BIT3 = "FALSE";
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [3:0] SRIOV_CAP_ENABLE = 4'h0;
    parameter TL2CFG_IF_PARITY_CHK = "TRUE";
    parameter [1:0] TL_COMPLETION_RAM_NUM_TLPS = 2'h0;
    parameter [1:0] TL_COMPLETION_RAM_SIZE = 2'h1;
    parameter [11:0] TL_CREDITS_CD = 12'h000;
    parameter [7:0] TL_CREDITS_CH = 8'h00;
    parameter [11:0] TL_CREDITS_NPD = 12'h004;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [11:0] TL_CREDITS_PD = 12'h0E0;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TIME = 5'h02;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT = 5'h08;
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter [0:0] TL_POSTED_RAM_SIZE = 1'h0;
    parameter TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TL_TX_TLP_STRADDLE_ENABLE = "FALSE";
    parameter TL_TX_TLP_TERMINATE_PARITY = "FALSE";
    parameter [15:0] TL_USER_SPARE = 16'h0000;
    parameter TPH_FROM_RAM_PIPELINE = "FALSE";
    parameter TPH_TO_RAM_PIPELINE = "FALSE";
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h80;
    parameter [11:0] VFG0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] VFG3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    output [7:0] AXIUSEROUT;
    output [7:0] CFGBUSNUMBER;
    output [1:0] CFGCURRENTSPEED;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXVECPENDINGSTATUS;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output [4:0] CFGLOCALERROROUT;
    output CFGLOCALERRORVALID;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [1:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [12:0] CFGMSIXRAMADDRESS;
    output CFGMSIXRAMREADENABLE;
    output [3:0] CFGMSIXRAMWRITEBYTEENABLE;
    output [35:0] CFGMSIXRAMWRITEDATA;
    output [2:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [1:0] CFGRXPMSTATE;
    output [11:0] CFGTPHRAMADDRESS;
    output CFGTPHRAMREADENABLE;
    output [3:0] CFGTPHRAMWRITEBYTEENABLE;
    output [35:0] CFGTPHRAMWRITEDATA;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [1:0] CFGTXPMSTATE;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [31:0] DBGCTRL0OUT;
    output [31:0] DBGCTRL1OUT;
    output [255:0] DBGDATA0OUT;
    output [255:0] DBGDATA1OUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [87:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [8:0] MIREPLAYRAMADDRESS0;
    output [8:0] MIREPLAYRAMADDRESS1;
    output MIREPLAYRAMREADENABLE0;
    output MIREPLAYRAMREADENABLE1;
    output [127:0] MIREPLAYRAMWRITEDATA0;
    output [127:0] MIREPLAYRAMWRITEDATA1;
    output MIREPLAYRAMWRITEENABLE0;
    output MIREPLAYRAMWRITEENABLE1;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS1;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE0;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE1;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS1;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA0;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA1;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE0;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS1;
    output MIRXPOSTEDREQUESTRAMREADENABLE0;
    output MIRXPOSTEDREQUESTRAMREADENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS1;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA0;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA1;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE0;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE1;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [5:0] PCIERQSEQNUM0;
    output [5:0] PCIERQSEQNUM1;
    output PCIERQSEQNUMVLD0;
    output PCIERQSEQNUMVLD1;
    output [7:0] PCIERQTAG0;
    output [7:0] PCIERQTAG1;
    output [3:0] PCIERQTAGAV;
    output PCIERQTAGVLD0;
    output PCIERQTAGVLD1;
    output [3:0] PCIETFCNPDAV;
    output [3:0] PCIETFCNPHAV;
    output [1:0] PIPERX00EQCONTROL;
    output PIPERX00POLARITY;
    output [1:0] PIPERX01EQCONTROL;
    output PIPERX01POLARITY;
    output [1:0] PIPERX02EQCONTROL;
    output PIPERX02POLARITY;
    output [1:0] PIPERX03EQCONTROL;
    output PIPERX03POLARITY;
    output [1:0] PIPERX04EQCONTROL;
    output PIPERX04POLARITY;
    output [1:0] PIPERX05EQCONTROL;
    output PIPERX05POLARITY;
    output [1:0] PIPERX06EQCONTROL;
    output PIPERX06POLARITY;
    output [1:0] PIPERX07EQCONTROL;
    output PIPERX07POLARITY;
    output [1:0] PIPERX08EQCONTROL;
    output PIPERX08POLARITY;
    output [1:0] PIPERX09EQCONTROL;
    output PIPERX09POLARITY;
    output [1:0] PIPERX10EQCONTROL;
    output PIPERX10POLARITY;
    output [1:0] PIPERX11EQCONTROL;
    output PIPERX11POLARITY;
    output [1:0] PIPERX12EQCONTROL;
    output PIPERX12POLARITY;
    output [1:0] PIPERX13EQCONTROL;
    output PIPERX13POLARITY;
    output [1:0] PIPERX14EQCONTROL;
    output PIPERX14POLARITY;
    output [1:0] PIPERX15EQCONTROL;
    output PIPERX15POLARITY;
    output [5:0] PIPERXEQLPLFFS;
    output [3:0] PIPERXEQLPTXPRESET;
    output [1:0] PIPETX00CHARISK;
    output PIPETX00COMPLIANCE;
    output [31:0] PIPETX00DATA;
    output PIPETX00DATAVALID;
    output PIPETX00ELECIDLE;
    output [1:0] PIPETX00EQCONTROL;
    output [5:0] PIPETX00EQDEEMPH;
    output [1:0] PIPETX00POWERDOWN;
    output PIPETX00STARTBLOCK;
    output [1:0] PIPETX00SYNCHEADER;
    output [1:0] PIPETX01CHARISK;
    output PIPETX01COMPLIANCE;
    output [31:0] PIPETX01DATA;
    output PIPETX01DATAVALID;
    output PIPETX01ELECIDLE;
    output [1:0] PIPETX01EQCONTROL;
    output [5:0] PIPETX01EQDEEMPH;
    output [1:0] PIPETX01POWERDOWN;
    output PIPETX01STARTBLOCK;
    output [1:0] PIPETX01SYNCHEADER;
    output [1:0] PIPETX02CHARISK;
    output PIPETX02COMPLIANCE;
    output [31:0] PIPETX02DATA;
    output PIPETX02DATAVALID;
    output PIPETX02ELECIDLE;
    output [1:0] PIPETX02EQCONTROL;
    output [5:0] PIPETX02EQDEEMPH;
    output [1:0] PIPETX02POWERDOWN;
    output PIPETX02STARTBLOCK;
    output [1:0] PIPETX02SYNCHEADER;
    output [1:0] PIPETX03CHARISK;
    output PIPETX03COMPLIANCE;
    output [31:0] PIPETX03DATA;
    output PIPETX03DATAVALID;
    output PIPETX03ELECIDLE;
    output [1:0] PIPETX03EQCONTROL;
    output [5:0] PIPETX03EQDEEMPH;
    output [1:0] PIPETX03POWERDOWN;
    output PIPETX03STARTBLOCK;
    output [1:0] PIPETX03SYNCHEADER;
    output [1:0] PIPETX04CHARISK;
    output PIPETX04COMPLIANCE;
    output [31:0] PIPETX04DATA;
    output PIPETX04DATAVALID;
    output PIPETX04ELECIDLE;
    output [1:0] PIPETX04EQCONTROL;
    output [5:0] PIPETX04EQDEEMPH;
    output [1:0] PIPETX04POWERDOWN;
    output PIPETX04STARTBLOCK;
    output [1:0] PIPETX04SYNCHEADER;
    output [1:0] PIPETX05CHARISK;
    output PIPETX05COMPLIANCE;
    output [31:0] PIPETX05DATA;
    output PIPETX05DATAVALID;
    output PIPETX05ELECIDLE;
    output [1:0] PIPETX05EQCONTROL;
    output [5:0] PIPETX05EQDEEMPH;
    output [1:0] PIPETX05POWERDOWN;
    output PIPETX05STARTBLOCK;
    output [1:0] PIPETX05SYNCHEADER;
    output [1:0] PIPETX06CHARISK;
    output PIPETX06COMPLIANCE;
    output [31:0] PIPETX06DATA;
    output PIPETX06DATAVALID;
    output PIPETX06ELECIDLE;
    output [1:0] PIPETX06EQCONTROL;
    output [5:0] PIPETX06EQDEEMPH;
    output [1:0] PIPETX06POWERDOWN;
    output PIPETX06STARTBLOCK;
    output [1:0] PIPETX06SYNCHEADER;
    output [1:0] PIPETX07CHARISK;
    output PIPETX07COMPLIANCE;
    output [31:0] PIPETX07DATA;
    output PIPETX07DATAVALID;
    output PIPETX07ELECIDLE;
    output [1:0] PIPETX07EQCONTROL;
    output [5:0] PIPETX07EQDEEMPH;
    output [1:0] PIPETX07POWERDOWN;
    output PIPETX07STARTBLOCK;
    output [1:0] PIPETX07SYNCHEADER;
    output [1:0] PIPETX08CHARISK;
    output PIPETX08COMPLIANCE;
    output [31:0] PIPETX08DATA;
    output PIPETX08DATAVALID;
    output PIPETX08ELECIDLE;
    output [1:0] PIPETX08EQCONTROL;
    output [5:0] PIPETX08EQDEEMPH;
    output [1:0] PIPETX08POWERDOWN;
    output PIPETX08STARTBLOCK;
    output [1:0] PIPETX08SYNCHEADER;
    output [1:0] PIPETX09CHARISK;
    output PIPETX09COMPLIANCE;
    output [31:0] PIPETX09DATA;
    output PIPETX09DATAVALID;
    output PIPETX09ELECIDLE;
    output [1:0] PIPETX09EQCONTROL;
    output [5:0] PIPETX09EQDEEMPH;
    output [1:0] PIPETX09POWERDOWN;
    output PIPETX09STARTBLOCK;
    output [1:0] PIPETX09SYNCHEADER;
    output [1:0] PIPETX10CHARISK;
    output PIPETX10COMPLIANCE;
    output [31:0] PIPETX10DATA;
    output PIPETX10DATAVALID;
    output PIPETX10ELECIDLE;
    output [1:0] PIPETX10EQCONTROL;
    output [5:0] PIPETX10EQDEEMPH;
    output [1:0] PIPETX10POWERDOWN;
    output PIPETX10STARTBLOCK;
    output [1:0] PIPETX10SYNCHEADER;
    output [1:0] PIPETX11CHARISK;
    output PIPETX11COMPLIANCE;
    output [31:0] PIPETX11DATA;
    output PIPETX11DATAVALID;
    output PIPETX11ELECIDLE;
    output [1:0] PIPETX11EQCONTROL;
    output [5:0] PIPETX11EQDEEMPH;
    output [1:0] PIPETX11POWERDOWN;
    output PIPETX11STARTBLOCK;
    output [1:0] PIPETX11SYNCHEADER;
    output [1:0] PIPETX12CHARISK;
    output PIPETX12COMPLIANCE;
    output [31:0] PIPETX12DATA;
    output PIPETX12DATAVALID;
    output PIPETX12ELECIDLE;
    output [1:0] PIPETX12EQCONTROL;
    output [5:0] PIPETX12EQDEEMPH;
    output [1:0] PIPETX12POWERDOWN;
    output PIPETX12STARTBLOCK;
    output [1:0] PIPETX12SYNCHEADER;
    output [1:0] PIPETX13CHARISK;
    output PIPETX13COMPLIANCE;
    output [31:0] PIPETX13DATA;
    output PIPETX13DATAVALID;
    output PIPETX13ELECIDLE;
    output [1:0] PIPETX13EQCONTROL;
    output [5:0] PIPETX13EQDEEMPH;
    output [1:0] PIPETX13POWERDOWN;
    output PIPETX13STARTBLOCK;
    output [1:0] PIPETX13SYNCHEADER;
    output [1:0] PIPETX14CHARISK;
    output PIPETX14COMPLIANCE;
    output [31:0] PIPETX14DATA;
    output PIPETX14DATAVALID;
    output PIPETX14ELECIDLE;
    output [1:0] PIPETX14EQCONTROL;
    output [5:0] PIPETX14EQDEEMPH;
    output [1:0] PIPETX14POWERDOWN;
    output PIPETX14STARTBLOCK;
    output [1:0] PIPETX14SYNCHEADER;
    output [1:0] PIPETX15CHARISK;
    output PIPETX15COMPLIANCE;
    output [31:0] PIPETX15DATA;
    output PIPETX15DATAVALID;
    output PIPETX15ELECIDLE;
    output [1:0] PIPETX15EQCONTROL;
    output [5:0] PIPETX15EQDEEMPH;
    output [1:0] PIPETX15POWERDOWN;
    output PIPETX15STARTBLOCK;
    output [1:0] PIPETX15SYNCHEADER;
    output PIPETXDEEMPH;
    output [2:0] PIPETXMARGIN;
    output [1:0] PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output PLGEN34EQMISMATCH;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [31:0] USERSPAREOUT;
    input [7:0] AXIUSERIN;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVIDPF0;
    input [15:0] CFGDEVIDPF1;
    input [15:0] CFGDEVIDPF2;
    input [15:0] CFGDEVIDPF3;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [7:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [1:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [1:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [7:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [1:0] CFGINTERRUPTMSIXVECPENDING;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [9:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTDEBUGACCESS;
    input [7:0] CFGMGMTFUNCTIONNUMBER;
    input CFGMGMTREAD;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [35:0] CFGMSIXRAMREADDATA;
    input CFGPMASPML1ENTRYREJECT;
    input CFGPMASPMTXL0SENTRYDISABLE;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVIDPF0;
    input [7:0] CFGREVIDPF1;
    input [7:0] CFGREVIDPF2;
    input [7:0] CFGREVIDPF3;
    input [15:0] CFGSUBSYSIDPF0;
    input [15:0] CFGSUBSYSIDPF1;
    input [15:0] CFGSUBSYSIDPF2;
    input [15:0] CFGSUBSYSIDPF3;
    input [15:0] CFGSUBSYSVENDID;
    input [35:0] CFGTPHRAMREADDATA;
    input [15:0] CFGVENDID;
    input CFGVFFLRDONE;
    input [7:0] CFGVFFLRFUNCNUM;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKMIREPLAYRAM0;
    input CORECLKMIREPLAYRAM1;
    input CORECLKMIRXCOMPLETIONRAM0;
    input CORECLKMIRXCOMPLETIONRAM1;
    input CORECLKMIRXPOSTEDREQUESTRAM0;
    input CORECLKMIRXPOSTEDREQUESTRAM1;
    input [5:0] DBGSEL0;
    input [5:0] DBGSEL1;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [5:0] MIREPLAYRAMERRCOR;
    input [5:0] MIREPLAYRAMERRUNCOR;
    input [127:0] MIREPLAYRAMREADDATA0;
    input [127:0] MIREPLAYRAMREADDATA1;
    input [11:0] MIRXCOMPLETIONRAMERRCOR;
    input [11:0] MIRXCOMPLETIONRAMERRUNCOR;
    input [143:0] MIRXCOMPLETIONRAMREADDATA0;
    input [143:0] MIRXCOMPLETIONRAMREADDATA1;
    input [5:0] MIRXPOSTEDREQUESTRAMERRCOR;
    input [5:0] MIRXPOSTEDREQUESTRAMERRUNCOR;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA0;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA1;
    input [1:0] PCIECOMPLDELIVERED;
    input [7:0] PCIECOMPLDELIVEREDTAG0;
    input [7:0] PCIECOMPLDELIVEREDTAG1;
    input [1:0] PCIECQNPREQ;
    input PCIECQNPUSERCREDITRCVD;
    input PCIECQPIPELINEEMPTY;
    input PCIEPOSTEDREQDELIVERED;
    input PIPECLK;
    input PIPECLKEN;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX00CHARISK;
    input [31:0] PIPERX00DATA;
    input PIPERX00DATAVALID;
    input PIPERX00ELECIDLE;
    input PIPERX00EQDONE;
    input PIPERX00EQLPADAPTDONE;
    input PIPERX00EQLPLFFSSEL;
    input [17:0] PIPERX00EQLPNEWTXCOEFFORPRESET;
    input PIPERX00PHYSTATUS;
    input [1:0] PIPERX00STARTBLOCK;
    input [2:0] PIPERX00STATUS;
    input [1:0] PIPERX00SYNCHEADER;
    input PIPERX00VALID;
    input [1:0] PIPERX01CHARISK;
    input [31:0] PIPERX01DATA;
    input PIPERX01DATAVALID;
    input PIPERX01ELECIDLE;
    input PIPERX01EQDONE;
    input PIPERX01EQLPADAPTDONE;
    input PIPERX01EQLPLFFSSEL;
    input [17:0] PIPERX01EQLPNEWTXCOEFFORPRESET;
    input PIPERX01PHYSTATUS;
    input [1:0] PIPERX01STARTBLOCK;
    input [2:0] PIPERX01STATUS;
    input [1:0] PIPERX01SYNCHEADER;
    input PIPERX01VALID;
    input [1:0] PIPERX02CHARISK;
    input [31:0] PIPERX02DATA;
    input PIPERX02DATAVALID;
    input PIPERX02ELECIDLE;
    input PIPERX02EQDONE;
    input PIPERX02EQLPADAPTDONE;
    input PIPERX02EQLPLFFSSEL;
    input [17:0] PIPERX02EQLPNEWTXCOEFFORPRESET;
    input PIPERX02PHYSTATUS;
    input [1:0] PIPERX02STARTBLOCK;
    input [2:0] PIPERX02STATUS;
    input [1:0] PIPERX02SYNCHEADER;
    input PIPERX02VALID;
    input [1:0] PIPERX03CHARISK;
    input [31:0] PIPERX03DATA;
    input PIPERX03DATAVALID;
    input PIPERX03ELECIDLE;
    input PIPERX03EQDONE;
    input PIPERX03EQLPADAPTDONE;
    input PIPERX03EQLPLFFSSEL;
    input [17:0] PIPERX03EQLPNEWTXCOEFFORPRESET;
    input PIPERX03PHYSTATUS;
    input [1:0] PIPERX03STARTBLOCK;
    input [2:0] PIPERX03STATUS;
    input [1:0] PIPERX03SYNCHEADER;
    input PIPERX03VALID;
    input [1:0] PIPERX04CHARISK;
    input [31:0] PIPERX04DATA;
    input PIPERX04DATAVALID;
    input PIPERX04ELECIDLE;
    input PIPERX04EQDONE;
    input PIPERX04EQLPADAPTDONE;
    input PIPERX04EQLPLFFSSEL;
    input [17:0] PIPERX04EQLPNEWTXCOEFFORPRESET;
    input PIPERX04PHYSTATUS;
    input [1:0] PIPERX04STARTBLOCK;
    input [2:0] PIPERX04STATUS;
    input [1:0] PIPERX04SYNCHEADER;
    input PIPERX04VALID;
    input [1:0] PIPERX05CHARISK;
    input [31:0] PIPERX05DATA;
    input PIPERX05DATAVALID;
    input PIPERX05ELECIDLE;
    input PIPERX05EQDONE;
    input PIPERX05EQLPADAPTDONE;
    input PIPERX05EQLPLFFSSEL;
    input [17:0] PIPERX05EQLPNEWTXCOEFFORPRESET;
    input PIPERX05PHYSTATUS;
    input [1:0] PIPERX05STARTBLOCK;
    input [2:0] PIPERX05STATUS;
    input [1:0] PIPERX05SYNCHEADER;
    input PIPERX05VALID;
    input [1:0] PIPERX06CHARISK;
    input [31:0] PIPERX06DATA;
    input PIPERX06DATAVALID;
    input PIPERX06ELECIDLE;
    input PIPERX06EQDONE;
    input PIPERX06EQLPADAPTDONE;
    input PIPERX06EQLPLFFSSEL;
    input [17:0] PIPERX06EQLPNEWTXCOEFFORPRESET;
    input PIPERX06PHYSTATUS;
    input [1:0] PIPERX06STARTBLOCK;
    input [2:0] PIPERX06STATUS;
    input [1:0] PIPERX06SYNCHEADER;
    input PIPERX06VALID;
    input [1:0] PIPERX07CHARISK;
    input [31:0] PIPERX07DATA;
    input PIPERX07DATAVALID;
    input PIPERX07ELECIDLE;
    input PIPERX07EQDONE;
    input PIPERX07EQLPADAPTDONE;
    input PIPERX07EQLPLFFSSEL;
    input [17:0] PIPERX07EQLPNEWTXCOEFFORPRESET;
    input PIPERX07PHYSTATUS;
    input [1:0] PIPERX07STARTBLOCK;
    input [2:0] PIPERX07STATUS;
    input [1:0] PIPERX07SYNCHEADER;
    input PIPERX07VALID;
    input [1:0] PIPERX08CHARISK;
    input [31:0] PIPERX08DATA;
    input PIPERX08DATAVALID;
    input PIPERX08ELECIDLE;
    input PIPERX08EQDONE;
    input PIPERX08EQLPADAPTDONE;
    input PIPERX08EQLPLFFSSEL;
    input [17:0] PIPERX08EQLPNEWTXCOEFFORPRESET;
    input PIPERX08PHYSTATUS;
    input [1:0] PIPERX08STARTBLOCK;
    input [2:0] PIPERX08STATUS;
    input [1:0] PIPERX08SYNCHEADER;
    input PIPERX08VALID;
    input [1:0] PIPERX09CHARISK;
    input [31:0] PIPERX09DATA;
    input PIPERX09DATAVALID;
    input PIPERX09ELECIDLE;
    input PIPERX09EQDONE;
    input PIPERX09EQLPADAPTDONE;
    input PIPERX09EQLPLFFSSEL;
    input [17:0] PIPERX09EQLPNEWTXCOEFFORPRESET;
    input PIPERX09PHYSTATUS;
    input [1:0] PIPERX09STARTBLOCK;
    input [2:0] PIPERX09STATUS;
    input [1:0] PIPERX09SYNCHEADER;
    input PIPERX09VALID;
    input [1:0] PIPERX10CHARISK;
    input [31:0] PIPERX10DATA;
    input PIPERX10DATAVALID;
    input PIPERX10ELECIDLE;
    input PIPERX10EQDONE;
    input PIPERX10EQLPADAPTDONE;
    input PIPERX10EQLPLFFSSEL;
    input [17:0] PIPERX10EQLPNEWTXCOEFFORPRESET;
    input PIPERX10PHYSTATUS;
    input [1:0] PIPERX10STARTBLOCK;
    input [2:0] PIPERX10STATUS;
    input [1:0] PIPERX10SYNCHEADER;
    input PIPERX10VALID;
    input [1:0] PIPERX11CHARISK;
    input [31:0] PIPERX11DATA;
    input PIPERX11DATAVALID;
    input PIPERX11ELECIDLE;
    input PIPERX11EQDONE;
    input PIPERX11EQLPADAPTDONE;
    input PIPERX11EQLPLFFSSEL;
    input [17:0] PIPERX11EQLPNEWTXCOEFFORPRESET;
    input PIPERX11PHYSTATUS;
    input [1:0] PIPERX11STARTBLOCK;
    input [2:0] PIPERX11STATUS;
    input [1:0] PIPERX11SYNCHEADER;
    input PIPERX11VALID;
    input [1:0] PIPERX12CHARISK;
    input [31:0] PIPERX12DATA;
    input PIPERX12DATAVALID;
    input PIPERX12ELECIDLE;
    input PIPERX12EQDONE;
    input PIPERX12EQLPADAPTDONE;
    input PIPERX12EQLPLFFSSEL;
    input [17:0] PIPERX12EQLPNEWTXCOEFFORPRESET;
    input PIPERX12PHYSTATUS;
    input [1:0] PIPERX12STARTBLOCK;
    input [2:0] PIPERX12STATUS;
    input [1:0] PIPERX12SYNCHEADER;
    input PIPERX12VALID;
    input [1:0] PIPERX13CHARISK;
    input [31:0] PIPERX13DATA;
    input PIPERX13DATAVALID;
    input PIPERX13ELECIDLE;
    input PIPERX13EQDONE;
    input PIPERX13EQLPADAPTDONE;
    input PIPERX13EQLPLFFSSEL;
    input [17:0] PIPERX13EQLPNEWTXCOEFFORPRESET;
    input PIPERX13PHYSTATUS;
    input [1:0] PIPERX13STARTBLOCK;
    input [2:0] PIPERX13STATUS;
    input [1:0] PIPERX13SYNCHEADER;
    input PIPERX13VALID;
    input [1:0] PIPERX14CHARISK;
    input [31:0] PIPERX14DATA;
    input PIPERX14DATAVALID;
    input PIPERX14ELECIDLE;
    input PIPERX14EQDONE;
    input PIPERX14EQLPADAPTDONE;
    input PIPERX14EQLPLFFSSEL;
    input [17:0] PIPERX14EQLPNEWTXCOEFFORPRESET;
    input PIPERX14PHYSTATUS;
    input [1:0] PIPERX14STARTBLOCK;
    input [2:0] PIPERX14STATUS;
    input [1:0] PIPERX14SYNCHEADER;
    input PIPERX14VALID;
    input [1:0] PIPERX15CHARISK;
    input [31:0] PIPERX15DATA;
    input PIPERX15DATAVALID;
    input PIPERX15ELECIDLE;
    input PIPERX15EQDONE;
    input PIPERX15EQLPADAPTDONE;
    input PIPERX15EQLPLFFSSEL;
    input [17:0] PIPERX15EQLPNEWTXCOEFFORPRESET;
    input PIPERX15PHYSTATUS;
    input [1:0] PIPERX15STARTBLOCK;
    input [2:0] PIPERX15STATUS;
    input [1:0] PIPERX15SYNCHEADER;
    input PIPERX15VALID;
    input [17:0] PIPETX00EQCOEFF;
    input PIPETX00EQDONE;
    input [17:0] PIPETX01EQCOEFF;
    input PIPETX01EQDONE;
    input [17:0] PIPETX02EQCOEFF;
    input PIPETX02EQDONE;
    input [17:0] PIPETX03EQCOEFF;
    input PIPETX03EQDONE;
    input [17:0] PIPETX04EQCOEFF;
    input PIPETX04EQDONE;
    input [17:0] PIPETX05EQCOEFF;
    input PIPETX05EQDONE;
    input [17:0] PIPETX06EQCOEFF;
    input PIPETX06EQDONE;
    input [17:0] PIPETX07EQCOEFF;
    input PIPETX07EQDONE;
    input [17:0] PIPETX08EQCOEFF;
    input PIPETX08EQDONE;
    input [17:0] PIPETX09EQCOEFF;
    input PIPETX09EQDONE;
    input [17:0] PIPETX10EQCOEFF;
    input PIPETX10EQDONE;
    input [17:0] PIPETX11EQCOEFF;
    input PIPETX11EQDONE;
    input [17:0] PIPETX12EQCOEFF;
    input PIPETX12EQDONE;
    input [17:0] PIPETX13EQCOEFF;
    input PIPETX13EQDONE;
    input [17:0] PIPETX14EQCOEFF;
    input PIPETX14EQDONE;
    input [17:0] PIPETX15EQCOEFF;
    input PIPETX15EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input PLGEN34REDOEQSPEED;
    input PLGEN34REDOEQUALIZATION;
    input RESETN;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [61:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input USERCLK;
    input USERCLK2;
    input USERCLKEN;
    input [31:0] USERSPAREIN;
endmodule

module PCIE4CE4 (...);
    parameter ARI_CAP_ENABLE = "FALSE";
    parameter AUTO_FLR_RESPONSE = "FALSE";
    parameter [7:0] AXISTEN_IF_CCIX_RX_CREDIT_LIMIT = 8'h08;
    parameter [7:0] AXISTEN_IF_CCIX_TX_CREDIT_LIMIT = 8'h08;
    parameter AXISTEN_IF_CCIX_TX_REGISTERED_TREADY = "FALSE";
    parameter [1:0] AXISTEN_IF_CC_ALIGNMENT_MODE = 2'h0;
    parameter [23:0] AXISTEN_IF_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
    parameter [27:0] AXISTEN_IF_COMPL_TIMEOUT_REG1 = 28'h2FAF080;
    parameter [1:0] AXISTEN_IF_CQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_CQ_EN_POISONED_MEM_WR = "FALSE";
    parameter AXISTEN_IF_ENABLE_256_TAGS = "FALSE";
    parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
    parameter AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE = "FALSE";
    parameter AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK = "TRUE";
    parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
    parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
    parameter AXISTEN_IF_EXT_512 = "FALSE";
    parameter AXISTEN_IF_EXT_512_CC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_CQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RC_STRADDLE = "FALSE";
    parameter AXISTEN_IF_EXT_512_RQ_STRADDLE = "FALSE";
    parameter AXISTEN_IF_LEGACY_MODE_ENABLE = "FALSE";
    parameter AXISTEN_IF_MSIX_FROM_RAM_PIPELINE = "FALSE";
    parameter AXISTEN_IF_MSIX_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_MSIX_TO_RAM_PIPELINE = "FALSE";
    parameter [1:0] AXISTEN_IF_RC_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
    parameter [1:0] AXISTEN_IF_RQ_ALIGNMENT_MODE = 2'h0;
    parameter AXISTEN_IF_RX_PARITY_EN = "TRUE";
    parameter AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT = "FALSE";
    parameter AXISTEN_IF_TX_PARITY_EN = "TRUE";
    parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
    parameter CCIX_DIRECT_ATTACH_MODE = "FALSE";
    parameter CCIX_ENABLE = "FALSE";
    parameter [15:0] CCIX_VENDOR_ID = 16'h0000;
    parameter CFG_BYPASS_MODE_ENABLE = "FALSE";
    parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
    parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
    parameter [15:0] DEBUG_AXI4ST_SPARE = 16'h0000;
    parameter [7:0] DEBUG_AXIST_DISABLE_FEATURE_BIT = 8'h00;
    parameter [3:0] DEBUG_CAR_SPARE = 4'h0;
    parameter [15:0] DEBUG_CFG_SPARE = 16'h0000;
    parameter [15:0] DEBUG_LL_SPARE = 16'h0000;
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL = "FALSE";
    parameter DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW = "FALSE";
    parameter DEBUG_PL_DISABLE_SCRAMBLING = "FALSE";
    parameter DEBUG_PL_SIM_RESET_LFSR = "FALSE";
    parameter [15:0] DEBUG_PL_SPARE = 16'h0000;
    parameter DEBUG_TL_DISABLE_FC_TIMEOUT = "FALSE";
    parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE";
    parameter [15:0] DEBUG_TL_SPARE = 16'h0000;
    parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
    parameter DSN_CAP_ENABLE = "FALSE";
    parameter EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter HEADER_TYPE_OVERRIDE = "FALSE";
    parameter IS_SWITCH_PORT = "FALSE";
    parameter LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
    parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
    parameter LL_ACK_TIMEOUT_EN = "FALSE";
    parameter integer LL_ACK_TIMEOUT_FUNC = 0;
    parameter LL_DISABLE_SCHED_TX_NAK = "FALSE";
    parameter LL_REPLAY_FROM_RAM_PIPELINE = "FALSE";
    parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
    parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
    parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
    parameter LL_REPLAY_TO_RAM_PIPELINE = "FALSE";
    parameter LL_RX_TLP_PARITY_GEN = "TRUE";
    parameter LL_TX_TLP_PARITY_CHK = "TRUE";
    parameter [15:0] LL_USER_SPARE = 16'h0000;
    parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h250;
    parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
    parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
    parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000;
    parameter MCAP_CONFIGURE_OVERRIDE = "FALSE";
    parameter MCAP_ENABLE = "FALSE";
    parameter MCAP_EOS_DESIGN_SWITCH = "FALSE";
    parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000;
    parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE";
    parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE";
    parameter [15:0] MCAP_VSEC_ID = 16'h0000;
    parameter [11:0] MCAP_VSEC_LEN = 12'h02C;
    parameter [3:0] MCAP_VSEC_REV = 4'h0;
    parameter PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE = "FALSE";
    parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
    parameter [4:0] PF0_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] PF0_ATS_CAP_NEXTPTR = 12'h000;
    parameter PF0_ATS_CAP_ON = "FALSE";
    parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF0_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF0_CLASS_CODE = 24'h000000;
    parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
    parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE";
    parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
    parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
    parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
    parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
    parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
    parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
    parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
    parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
    parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
    parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
    parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4 = 7;
    parameter [0:0] PF0_LINK_CONTROL_RCB = 1'h0;
    parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
    parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
    parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
    parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
    parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [5:0] PF0_MSIX_VECTOR_COUNT = 6'h04;
    parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF0_PM_CAP_ID = 8'h01;
    parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
    parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
    parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
    parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
    parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
    parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
    parameter [11:0] PF0_PRI_CAP_NEXTPTR = 12'h000;
    parameter PF0_PRI_CAP_ON = "FALSE";
    parameter [31:0] PF0_PRI_OST_PR_CAPACITY = 32'h00000000;
    parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000;
    parameter PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
    parameter PF0_TPHR_CAP_ENABLE = "FALSE";
    parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
    parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
    parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
    parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
    parameter [3:0] PF0_VC_ARB_CAPABILITY = 4'h0;
    parameter [7:0] PF0_VC_ARB_TBL_OFFSET = 8'h00;
    parameter PF0_VC_CAP_ENABLE = "FALSE";
    parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
    parameter [3:0] PF0_VC_CAP_VER = 4'h1;
    parameter PF0_VC_EXTENDED_COUNT = "FALSE";
    parameter PF0_VC_LOW_PRIORITY_EXTENDED_COUNT = "FALSE";
    parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [4:0] PF1_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] PF1_ATS_CAP_NEXTPTR = 12'h000;
    parameter PF1_ATS_CAP_ON = "FALSE";
    parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF1_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF1_CLASS_CODE = 24'h000000;
    parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF1_PRI_CAP_NEXTPTR = 12'h000;
    parameter PF1_PRI_CAP_ON = "FALSE";
    parameter [31:0] PF1_PRI_OST_PR_CAPACITY = 32'h00000000;
    parameter PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [4:0] PF2_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] PF2_ATS_CAP_NEXTPTR = 12'h000;
    parameter PF2_ATS_CAP_ON = "FALSE";
    parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF2_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF2_CLASS_CODE = 24'h000000;
    parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF2_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF2_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF2_PRI_CAP_NEXTPTR = 12'h000;
    parameter PF2_PRI_CAP_ON = "FALSE";
    parameter [31:0] PF2_PRI_OST_PR_CAPACITY = 32'h00000000;
    parameter PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000;
    parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00;
    parameter [4:0] PF3_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] PF3_ATS_CAP_NEXTPTR = 12'h000;
    parameter PF3_ATS_CAP_ON = "FALSE";
    parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_BAR5_CONTROL = 3'h0;
    parameter [7:0] PF3_CAPABILITY_POINTER = 8'h80;
    parameter [23:0] PF3_CLASS_CODE = 24'h000000;
    parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
    parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C;
    parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
    parameter PF3_EXPANSION_ROM_ENABLE = "FALSE";
    parameter [2:0] PF3_INTERRUPT_PIN = 3'h1;
    parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer PF3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer PF3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0;
    parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00;
    parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE";
    parameter [7:0] PF3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00;
    parameter [11:0] PF3_PRI_CAP_NEXTPTR = 12'h000;
    parameter PF3_PRI_CAP_ON = "FALSE";
    parameter [31:0] PF3_PRI_OST_PR_CAPACITY = 32'h00000000;
    parameter PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED = "FALSE";
    parameter [5:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
    parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0;
    parameter [5:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 6'h03;
    parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4;
    parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
    parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0;
    parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000;
    parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000;
    parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000;
    parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1;
    parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000;
    parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000;
    parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
    parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000;
    parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter PL_CFG_STATE_ROBUSTNESS_ENABLE = "TRUE";
    parameter PL_CTRL_SKP_GEN_ENABLE = "FALSE";
    parameter PL_CTRL_SKP_PARITY_AND_CRC_CHECK_DISABLE = "TRUE";
    parameter PL_DEEMPH_SOURCE_SELECT = "TRUE";
    parameter PL_DESKEW_ON_SKIP_IN_GEN12 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE";
    parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4 = "FALSE";
    parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE";
    parameter PL_DISABLE_DC_BALANCE = "FALSE";
    parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
    parameter PL_DISABLE_LANE_REVERSAL = "FALSE";
    parameter [1:0] PL_DISABLE_LFSR_UPDATE_ON_SKP = 2'h0;
    parameter PL_DISABLE_RETRAIN_ON_EB_ERROR = "FALSE";
    parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE";
    parameter [15:0] PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR = 16'h0000;
    parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
    parameter [1:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK = 2'h0;
    parameter [1:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK = 2'h0;
    parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
    parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
    parameter [1:0] PL_EQ_BYPASS_PHASE23 = 2'h0;
    parameter [5:0] PL_EQ_DEFAULT_RX_PRESET_HINT = 6'h33;
    parameter [7:0] PL_EQ_DEFAULT_TX_PRESET = 8'h44;
    parameter PL_EQ_DISABLE_MISMATCH_CHECK = "TRUE";
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE0 = 2'h0;
    parameter [1:0] PL_EQ_RX_ADAPT_EQ_PHASE1 = 2'h0;
    parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
    parameter PL_EQ_TX_8G_EQ_TS2_ENABLE = "FALSE";
    parameter PL_EXIT_LOOPBACK_ON_EI_ENTRY = "TRUE";
    parameter PL_INFER_EI_DISABLE_LPBK_ACTIVE = "TRUE";
    parameter PL_INFER_EI_DISABLE_REC_RC = "FALSE";
    parameter PL_INFER_EI_DISABLE_REC_SPD = "FALSE";
    parameter [31:0] PL_LANE0_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE10_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE11_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE12_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE13_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE14_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE15_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE1_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE2_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE3_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE4_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE5_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE6_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE7_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE8_EQ_CONTROL = 32'h00003F00;
    parameter [31:0] PL_LANE9_EQ_CONTROL = 32'h00003F00;
    parameter [3:0] PL_LINK_CAP_MAX_LINK_SPEED = 4'h4;
    parameter [4:0] PL_LINK_CAP_MAX_LINK_WIDTH = 5'h08;
    parameter integer PL_N_FTS = 255;
    parameter PL_QUIESCE_GUARANTEE_DISABLE = "FALSE";
    parameter PL_REDO_EQ_SOURCE_SELECT = "TRUE";
    parameter [7:0] PL_REPORT_ALL_PHY_ERRORS = 8'h00;
    parameter [1:0] PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_CLWS_GEN4 = 4'h0;
    parameter [1:0] PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS = 2'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN3 = 4'h0;
    parameter [3:0] PL_RX_ADAPT_TIMER_RRL_GEN4 = 4'h0;
    parameter [1:0] PL_RX_L0S_EXIT_TO_RECOVERY = 2'h0;
    parameter [1:0] PL_SIM_FAST_LINK_TRAINING = 2'h0;
    parameter PL_SRIS_ENABLE = "FALSE";
    parameter [6:0] PL_SRIS_SKPOS_GEN_SPD_VEC = 7'h00;
    parameter [6:0] PL_SRIS_SKPOS_REC_SPD_VEC = 7'h00;
    parameter PL_UPSTREAM_FACING = "TRUE";
    parameter [15:0] PL_USER_SPARE = 16'h0000;
    parameter [15:0] PL_USER_SPARE2 = 16'h0000;
    parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h1500;
    parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h003E8;
    parameter PM_ENABLE_L23_ENTRY = "FALSE";
    parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
    parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000100;
    parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h00000;
    parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0100;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000;
    parameter SIM_VERSION = "1.0";
    parameter SPARE_BIT0 = "FALSE";
    parameter integer SPARE_BIT1 = 0;
    parameter integer SPARE_BIT2 = 0;
    parameter SPARE_BIT3 = "FALSE";
    parameter integer SPARE_BIT4 = 0;
    parameter integer SPARE_BIT5 = 0;
    parameter integer SPARE_BIT6 = 0;
    parameter integer SPARE_BIT7 = 0;
    parameter integer SPARE_BIT8 = 0;
    parameter [7:0] SPARE_BYTE0 = 8'h00;
    parameter [7:0] SPARE_BYTE1 = 8'h00;
    parameter [7:0] SPARE_BYTE2 = 8'h00;
    parameter [7:0] SPARE_BYTE3 = 8'h00;
    parameter [31:0] SPARE_WORD0 = 32'h00000000;
    parameter [31:0] SPARE_WORD1 = 32'h00000000;
    parameter [31:0] SPARE_WORD2 = 32'h00000000;
    parameter [31:0] SPARE_WORD3 = 32'h00000000;
    parameter [3:0] SRIOV_CAP_ENABLE = 4'h0;
    parameter TL2CFG_IF_PARITY_CHK = "TRUE";
    parameter [1:0] TL_COMPLETION_RAM_NUM_TLPS = 2'h0;
    parameter [1:0] TL_COMPLETION_RAM_SIZE = 2'h1;
    parameter [11:0] TL_CREDITS_CD = 12'h000;
    parameter [11:0] TL_CREDITS_CD_VC1 = 12'h000;
    parameter [7:0] TL_CREDITS_CH = 8'h00;
    parameter [7:0] TL_CREDITS_CH_VC1 = 8'h00;
    parameter [11:0] TL_CREDITS_NPD = 12'h004;
    parameter [11:0] TL_CREDITS_NPD_VC1 = 12'h000;
    parameter [7:0] TL_CREDITS_NPH = 8'h20;
    parameter [7:0] TL_CREDITS_NPH_VC1 = 8'h01;
    parameter [11:0] TL_CREDITS_PD = 12'h0E0;
    parameter [11:0] TL_CREDITS_PD_VC1 = 12'h3E0;
    parameter [7:0] TL_CREDITS_PH = 8'h20;
    parameter [7:0] TL_CREDITS_PH_VC1 = 8'h20;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TIME = 5'h02;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TIME_VC1 = 5'h02;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT = 5'h08;
    parameter [4:0] TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT_VC1 = 5'h08;
    parameter TL_FEATURE_ENABLE_FC_SCALING = "FALSE";
    parameter [1:0] TL_PF_ENABLE_REG = 2'h0;
    parameter [0:0] TL_POSTED_RAM_SIZE = 1'h0;
    parameter TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_FROM_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_READ_PIPELINE = "FALSE";
    parameter TL_RX_POSTED_TO_RAM_WRITE_PIPELINE = "FALSE";
    parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE";
    parameter TL_TX_TLP_STRADDLE_ENABLE = "FALSE";
    parameter TL_TX_TLP_TERMINATE_PARITY = "FALSE";
    parameter [15:0] TL_USER_SPARE = 16'h0000;
    parameter TPH_FROM_RAM_PIPELINE = "FALSE";
    parameter TPH_TO_RAM_PIPELINE = "FALSE";
    parameter [7:0] VF0_CAPABILITY_POINTER = 8'h80;
    parameter [11:0] VFG0_ARI_CAP_NEXTPTR = 12'h000;
    parameter [4:0] VFG0_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] VFG0_ATS_CAP_NEXTPTR = 12'h000;
    parameter VFG0_ATS_CAP_ON = "FALSE";
    parameter [7:0] VFG0_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG0_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG0_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG0_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG0_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG0_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG0_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG1_ARI_CAP_NEXTPTR = 12'h000;
    parameter [4:0] VFG1_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] VFG1_ATS_CAP_NEXTPTR = 12'h000;
    parameter VFG1_ATS_CAP_ON = "FALSE";
    parameter [7:0] VFG1_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG1_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG1_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG1_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG1_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG1_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG1_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG2_ARI_CAP_NEXTPTR = 12'h000;
    parameter [4:0] VFG2_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] VFG2_ATS_CAP_NEXTPTR = 12'h000;
    parameter VFG2_ATS_CAP_ON = "FALSE";
    parameter [7:0] VFG2_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG2_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG2_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG2_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG2_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG2_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG2_TPHR_CAP_ST_MODE_SEL = 3'h0;
    parameter [11:0] VFG3_ARI_CAP_NEXTPTR = 12'h000;
    parameter [4:0] VFG3_ATS_CAP_INV_QUEUE_DEPTH = 5'h00;
    parameter [11:0] VFG3_ATS_CAP_NEXTPTR = 12'h000;
    parameter VFG3_ATS_CAP_ON = "FALSE";
    parameter [7:0] VFG3_MSIX_CAP_NEXTPTR = 8'h00;
    parameter integer VFG3_MSIX_CAP_PBA_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
    parameter integer VFG3_MSIX_CAP_TABLE_BIR = 0;
    parameter [28:0] VFG3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
    parameter [10:0] VFG3_MSIX_CAP_TABLE_SIZE = 11'h000;
    parameter [7:0] VFG3_PCIE_CAP_NEXTPTR = 8'h00;
    parameter [11:0] VFG3_TPHR_CAP_NEXTPTR = 12'h000;
    parameter [2:0] VFG3_TPHR_CAP_ST_MODE_SEL = 3'h0;
    output [7:0] AXIUSEROUT;
    output CCIXTXCREDIT;
    output [7:0] CFGBUSNUMBER;
    output [1:0] CFGCURRENTSPEED;
    output CFGERRCOROUT;
    output CFGERRFATALOUT;
    output CFGERRNONFATALOUT;
    output [7:0] CFGEXTFUNCTIONNUMBER;
    output CFGEXTREADRECEIVED;
    output [9:0] CFGEXTREGISTERNUMBER;
    output [3:0] CFGEXTWRITEBYTEENABLE;
    output [31:0] CFGEXTWRITEDATA;
    output CFGEXTWRITERECEIVED;
    output [11:0] CFGFCCPLD;
    output [7:0] CFGFCCPLH;
    output [11:0] CFGFCNPD;
    output [7:0] CFGFCNPH;
    output [11:0] CFGFCPD;
    output [7:0] CFGFCPH;
    output [3:0] CFGFLRINPROCESS;
    output [11:0] CFGFUNCTIONPOWERSTATE;
    output [15:0] CFGFUNCTIONSTATUS;
    output CFGHOTRESETOUT;
    output [31:0] CFGINTERRUPTMSIDATA;
    output [3:0] CFGINTERRUPTMSIENABLE;
    output CFGINTERRUPTMSIFAIL;
    output CFGINTERRUPTMSIMASKUPDATE;
    output [11:0] CFGINTERRUPTMSIMMENABLE;
    output CFGINTERRUPTMSISENT;
    output [3:0] CFGINTERRUPTMSIXENABLE;
    output [3:0] CFGINTERRUPTMSIXMASK;
    output CFGINTERRUPTMSIXVECPENDINGSTATUS;
    output CFGINTERRUPTSENT;
    output [1:0] CFGLINKPOWERSTATE;
    output [4:0] CFGLOCALERROROUT;
    output CFGLOCALERRORVALID;
    output CFGLTRENABLE;
    output [5:0] CFGLTSSMSTATE;
    output [1:0] CFGMAXPAYLOAD;
    output [2:0] CFGMAXREADREQ;
    output [31:0] CFGMGMTREADDATA;
    output CFGMGMTREADWRITEDONE;
    output CFGMSGRECEIVED;
    output [7:0] CFGMSGRECEIVEDDATA;
    output [4:0] CFGMSGRECEIVEDTYPE;
    output CFGMSGTRANSMITDONE;
    output [12:0] CFGMSIXRAMADDRESS;
    output CFGMSIXRAMREADENABLE;
    output [3:0] CFGMSIXRAMWRITEBYTEENABLE;
    output [35:0] CFGMSIXRAMWRITEDATA;
    output [2:0] CFGNEGOTIATEDWIDTH;
    output [1:0] CFGOBFFENABLE;
    output CFGPHYLINKDOWN;
    output [1:0] CFGPHYLINKSTATUS;
    output CFGPLSTATUSCHANGE;
    output CFGPOWERSTATECHANGEINTERRUPT;
    output [3:0] CFGRCBSTATUS;
    output [1:0] CFGRXPMSTATE;
    output [11:0] CFGTPHRAMADDRESS;
    output CFGTPHRAMREADENABLE;
    output [3:0] CFGTPHRAMWRITEBYTEENABLE;
    output [35:0] CFGTPHRAMWRITEDATA;
    output [3:0] CFGTPHREQUESTERENABLE;
    output [11:0] CFGTPHSTMODE;
    output [1:0] CFGTXPMSTATE;
    output CFGVC1ENABLE;
    output CFGVC1NEGOTIATIONPENDING;
    output CONFMCAPDESIGNSWITCH;
    output CONFMCAPEOS;
    output CONFMCAPINUSEBYPCIE;
    output CONFREQREADY;
    output [31:0] CONFRESPRDATA;
    output CONFRESPVALID;
    output [129:0] DBGCCIXOUT;
    output [31:0] DBGCTRL0OUT;
    output [31:0] DBGCTRL1OUT;
    output [255:0] DBGDATA0OUT;
    output [255:0] DBGDATA1OUT;
    output [15:0] DRPDO;
    output DRPRDY;
    output [45:0] MAXISCCIXRXTUSER;
    output MAXISCCIXRXTVALID;
    output [255:0] MAXISCQTDATA;
    output [7:0] MAXISCQTKEEP;
    output MAXISCQTLAST;
    output [87:0] MAXISCQTUSER;
    output MAXISCQTVALID;
    output [255:0] MAXISRCTDATA;
    output [7:0] MAXISRCTKEEP;
    output MAXISRCTLAST;
    output [74:0] MAXISRCTUSER;
    output MAXISRCTVALID;
    output [8:0] MIREPLAYRAMADDRESS0;
    output [8:0] MIREPLAYRAMADDRESS1;
    output MIREPLAYRAMREADENABLE0;
    output MIREPLAYRAMREADENABLE1;
    output [127:0] MIREPLAYRAMWRITEDATA0;
    output [127:0] MIREPLAYRAMWRITEDATA1;
    output MIREPLAYRAMWRITEENABLE0;
    output MIREPLAYRAMWRITEENABLE1;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMREADADDRESS1;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE0;
    output [1:0] MIRXCOMPLETIONRAMREADENABLE1;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS0;
    output [8:0] MIRXCOMPLETIONRAMWRITEADDRESS1;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA0;
    output [143:0] MIRXCOMPLETIONRAMWRITEDATA1;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE0;
    output [1:0] MIRXCOMPLETIONRAMWRITEENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMREADADDRESS1;
    output MIRXPOSTEDREQUESTRAMREADENABLE0;
    output MIRXPOSTEDREQUESTRAMREADENABLE1;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS0;
    output [8:0] MIRXPOSTEDREQUESTRAMWRITEADDRESS1;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA0;
    output [143:0] MIRXPOSTEDREQUESTRAMWRITEDATA1;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE0;
    output MIRXPOSTEDREQUESTRAMWRITEENABLE1;
    output [5:0] PCIECQNPREQCOUNT;
    output PCIEPERST0B;
    output PCIEPERST1B;
    output [5:0] PCIERQSEQNUM0;
    output [5:0] PCIERQSEQNUM1;
    output PCIERQSEQNUMVLD0;
    output PCIERQSEQNUMVLD1;
    output [7:0] PCIERQTAG0;
    output [7:0] PCIERQTAG1;
    output [3:0] PCIERQTAGAV;
    output PCIERQTAGVLD0;
    output PCIERQTAGVLD1;
    output [3:0] PCIETFCNPDAV;
    output [3:0] PCIETFCNPHAV;
    output [1:0] PIPERX00EQCONTROL;
    output PIPERX00POLARITY;
    output [1:0] PIPERX01EQCONTROL;
    output PIPERX01POLARITY;
    output [1:0] PIPERX02EQCONTROL;
    output PIPERX02POLARITY;
    output [1:0] PIPERX03EQCONTROL;
    output PIPERX03POLARITY;
    output [1:0] PIPERX04EQCONTROL;
    output PIPERX04POLARITY;
    output [1:0] PIPERX05EQCONTROL;
    output PIPERX05POLARITY;
    output [1:0] PIPERX06EQCONTROL;
    output PIPERX06POLARITY;
    output [1:0] PIPERX07EQCONTROL;
    output PIPERX07POLARITY;
    output [1:0] PIPERX08EQCONTROL;
    output PIPERX08POLARITY;
    output [1:0] PIPERX09EQCONTROL;
    output PIPERX09POLARITY;
    output [1:0] PIPERX10EQCONTROL;
    output PIPERX10POLARITY;
    output [1:0] PIPERX11EQCONTROL;
    output PIPERX11POLARITY;
    output [1:0] PIPERX12EQCONTROL;
    output PIPERX12POLARITY;
    output [1:0] PIPERX13EQCONTROL;
    output PIPERX13POLARITY;
    output [1:0] PIPERX14EQCONTROL;
    output PIPERX14POLARITY;
    output [1:0] PIPERX15EQCONTROL;
    output PIPERX15POLARITY;
    output [5:0] PIPERXEQLPLFFS;
    output [3:0] PIPERXEQLPTXPRESET;
    output [1:0] PIPETX00CHARISK;
    output PIPETX00COMPLIANCE;
    output [31:0] PIPETX00DATA;
    output PIPETX00DATAVALID;
    output PIPETX00ELECIDLE;
    output [1:0] PIPETX00EQCONTROL;
    output [5:0] PIPETX00EQDEEMPH;
    output [1:0] PIPETX00POWERDOWN;
    output PIPETX00STARTBLOCK;
    output [1:0] PIPETX00SYNCHEADER;
    output [1:0] PIPETX01CHARISK;
    output PIPETX01COMPLIANCE;
    output [31:0] PIPETX01DATA;
    output PIPETX01DATAVALID;
    output PIPETX01ELECIDLE;
    output [1:0] PIPETX01EQCONTROL;
    output [5:0] PIPETX01EQDEEMPH;
    output [1:0] PIPETX01POWERDOWN;
    output PIPETX01STARTBLOCK;
    output [1:0] PIPETX01SYNCHEADER;
    output [1:0] PIPETX02CHARISK;
    output PIPETX02COMPLIANCE;
    output [31:0] PIPETX02DATA;
    output PIPETX02DATAVALID;
    output PIPETX02ELECIDLE;
    output [1:0] PIPETX02EQCONTROL;
    output [5:0] PIPETX02EQDEEMPH;
    output [1:0] PIPETX02POWERDOWN;
    output PIPETX02STARTBLOCK;
    output [1:0] PIPETX02SYNCHEADER;
    output [1:0] PIPETX03CHARISK;
    output PIPETX03COMPLIANCE;
    output [31:0] PIPETX03DATA;
    output PIPETX03DATAVALID;
    output PIPETX03ELECIDLE;
    output [1:0] PIPETX03EQCONTROL;
    output [5:0] PIPETX03EQDEEMPH;
    output [1:0] PIPETX03POWERDOWN;
    output PIPETX03STARTBLOCK;
    output [1:0] PIPETX03SYNCHEADER;
    output [1:0] PIPETX04CHARISK;
    output PIPETX04COMPLIANCE;
    output [31:0] PIPETX04DATA;
    output PIPETX04DATAVALID;
    output PIPETX04ELECIDLE;
    output [1:0] PIPETX04EQCONTROL;
    output [5:0] PIPETX04EQDEEMPH;
    output [1:0] PIPETX04POWERDOWN;
    output PIPETX04STARTBLOCK;
    output [1:0] PIPETX04SYNCHEADER;
    output [1:0] PIPETX05CHARISK;
    output PIPETX05COMPLIANCE;
    output [31:0] PIPETX05DATA;
    output PIPETX05DATAVALID;
    output PIPETX05ELECIDLE;
    output [1:0] PIPETX05EQCONTROL;
    output [5:0] PIPETX05EQDEEMPH;
    output [1:0] PIPETX05POWERDOWN;
    output PIPETX05STARTBLOCK;
    output [1:0] PIPETX05SYNCHEADER;
    output [1:0] PIPETX06CHARISK;
    output PIPETX06COMPLIANCE;
    output [31:0] PIPETX06DATA;
    output PIPETX06DATAVALID;
    output PIPETX06ELECIDLE;
    output [1:0] PIPETX06EQCONTROL;
    output [5:0] PIPETX06EQDEEMPH;
    output [1:0] PIPETX06POWERDOWN;
    output PIPETX06STARTBLOCK;
    output [1:0] PIPETX06SYNCHEADER;
    output [1:0] PIPETX07CHARISK;
    output PIPETX07COMPLIANCE;
    output [31:0] PIPETX07DATA;
    output PIPETX07DATAVALID;
    output PIPETX07ELECIDLE;
    output [1:0] PIPETX07EQCONTROL;
    output [5:0] PIPETX07EQDEEMPH;
    output [1:0] PIPETX07POWERDOWN;
    output PIPETX07STARTBLOCK;
    output [1:0] PIPETX07SYNCHEADER;
    output [1:0] PIPETX08CHARISK;
    output PIPETX08COMPLIANCE;
    output [31:0] PIPETX08DATA;
    output PIPETX08DATAVALID;
    output PIPETX08ELECIDLE;
    output [1:0] PIPETX08EQCONTROL;
    output [5:0] PIPETX08EQDEEMPH;
    output [1:0] PIPETX08POWERDOWN;
    output PIPETX08STARTBLOCK;
    output [1:0] PIPETX08SYNCHEADER;
    output [1:0] PIPETX09CHARISK;
    output PIPETX09COMPLIANCE;
    output [31:0] PIPETX09DATA;
    output PIPETX09DATAVALID;
    output PIPETX09ELECIDLE;
    output [1:0] PIPETX09EQCONTROL;
    output [5:0] PIPETX09EQDEEMPH;
    output [1:0] PIPETX09POWERDOWN;
    output PIPETX09STARTBLOCK;
    output [1:0] PIPETX09SYNCHEADER;
    output [1:0] PIPETX10CHARISK;
    output PIPETX10COMPLIANCE;
    output [31:0] PIPETX10DATA;
    output PIPETX10DATAVALID;
    output PIPETX10ELECIDLE;
    output [1:0] PIPETX10EQCONTROL;
    output [5:0] PIPETX10EQDEEMPH;
    output [1:0] PIPETX10POWERDOWN;
    output PIPETX10STARTBLOCK;
    output [1:0] PIPETX10SYNCHEADER;
    output [1:0] PIPETX11CHARISK;
    output PIPETX11COMPLIANCE;
    output [31:0] PIPETX11DATA;
    output PIPETX11DATAVALID;
    output PIPETX11ELECIDLE;
    output [1:0] PIPETX11EQCONTROL;
    output [5:0] PIPETX11EQDEEMPH;
    output [1:0] PIPETX11POWERDOWN;
    output PIPETX11STARTBLOCK;
    output [1:0] PIPETX11SYNCHEADER;
    output [1:0] PIPETX12CHARISK;
    output PIPETX12COMPLIANCE;
    output [31:0] PIPETX12DATA;
    output PIPETX12DATAVALID;
    output PIPETX12ELECIDLE;
    output [1:0] PIPETX12EQCONTROL;
    output [5:0] PIPETX12EQDEEMPH;
    output [1:0] PIPETX12POWERDOWN;
    output PIPETX12STARTBLOCK;
    output [1:0] PIPETX12SYNCHEADER;
    output [1:0] PIPETX13CHARISK;
    output PIPETX13COMPLIANCE;
    output [31:0] PIPETX13DATA;
    output PIPETX13DATAVALID;
    output PIPETX13ELECIDLE;
    output [1:0] PIPETX13EQCONTROL;
    output [5:0] PIPETX13EQDEEMPH;
    output [1:0] PIPETX13POWERDOWN;
    output PIPETX13STARTBLOCK;
    output [1:0] PIPETX13SYNCHEADER;
    output [1:0] PIPETX14CHARISK;
    output PIPETX14COMPLIANCE;
    output [31:0] PIPETX14DATA;
    output PIPETX14DATAVALID;
    output PIPETX14ELECIDLE;
    output [1:0] PIPETX14EQCONTROL;
    output [5:0] PIPETX14EQDEEMPH;
    output [1:0] PIPETX14POWERDOWN;
    output PIPETX14STARTBLOCK;
    output [1:0] PIPETX14SYNCHEADER;
    output [1:0] PIPETX15CHARISK;
    output PIPETX15COMPLIANCE;
    output [31:0] PIPETX15DATA;
    output PIPETX15DATAVALID;
    output PIPETX15ELECIDLE;
    output [1:0] PIPETX15EQCONTROL;
    output [5:0] PIPETX15EQDEEMPH;
    output [1:0] PIPETX15POWERDOWN;
    output PIPETX15STARTBLOCK;
    output [1:0] PIPETX15SYNCHEADER;
    output PIPETXDEEMPH;
    output [2:0] PIPETXMARGIN;
    output [1:0] PIPETXRATE;
    output PIPETXRCVRDET;
    output PIPETXRESET;
    output PIPETXSWING;
    output PLEQINPROGRESS;
    output [1:0] PLEQPHASE;
    output PLGEN34EQMISMATCH;
    output [3:0] SAXISCCTREADY;
    output [3:0] SAXISRQTREADY;
    output [23:0] USERSPAREOUT;
    input [7:0] AXIUSERIN;
    input CCIXOPTIMIZEDTLPTXANDRXENABLE;
    input CCIXRXCORRECTABLEERRORDETECTED;
    input CCIXRXFIFOOVERFLOW;
    input CCIXRXTLPFORWARDED0;
    input CCIXRXTLPFORWARDED1;
    input [5:0] CCIXRXTLPFORWARDEDLENGTH0;
    input [5:0] CCIXRXTLPFORWARDEDLENGTH1;
    input CCIXRXUNCORRECTABLEERRORDETECTED;
    input CFGCONFIGSPACEENABLE;
    input [15:0] CFGDEVIDPF0;
    input [15:0] CFGDEVIDPF1;
    input [15:0] CFGDEVIDPF2;
    input [15:0] CFGDEVIDPF3;
    input [7:0] CFGDSBUSNUMBER;
    input [4:0] CFGDSDEVICENUMBER;
    input [2:0] CFGDSFUNCTIONNUMBER;
    input [63:0] CFGDSN;
    input [7:0] CFGDSPORTNUMBER;
    input CFGERRCORIN;
    input CFGERRUNCORIN;
    input [31:0] CFGEXTREADDATA;
    input CFGEXTREADDATAVALID;
    input [2:0] CFGFCSEL;
    input CFGFCVCSEL;
    input [3:0] CFGFLRDONE;
    input CFGHOTRESETIN;
    input [3:0] CFGINTERRUPTINT;
    input [2:0] CFGINTERRUPTMSIATTR;
    input [7:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
    input [31:0] CFGINTERRUPTMSIINT;
    input [31:0] CFGINTERRUPTMSIPENDINGSTATUS;
    input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
    input [1:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
    input [1:0] CFGINTERRUPTMSISELECT;
    input CFGINTERRUPTMSITPHPRESENT;
    input [7:0] CFGINTERRUPTMSITPHSTTAG;
    input [1:0] CFGINTERRUPTMSITPHTYPE;
    input [63:0] CFGINTERRUPTMSIXADDRESS;
    input [31:0] CFGINTERRUPTMSIXDATA;
    input CFGINTERRUPTMSIXINT;
    input [1:0] CFGINTERRUPTMSIXVECPENDING;
    input [3:0] CFGINTERRUPTPENDING;
    input CFGLINKTRAININGENABLE;
    input [9:0] CFGMGMTADDR;
    input [3:0] CFGMGMTBYTEENABLE;
    input CFGMGMTDEBUGACCESS;
    input [7:0] CFGMGMTFUNCTIONNUMBER;
    input CFGMGMTREAD;
    input CFGMGMTWRITE;
    input [31:0] CFGMGMTWRITEDATA;
    input CFGMSGTRANSMIT;
    input [31:0] CFGMSGTRANSMITDATA;
    input [2:0] CFGMSGTRANSMITTYPE;
    input [35:0] CFGMSIXRAMREADDATA;
    input CFGPMASPML1ENTRYREJECT;
    input CFGPMASPMTXL0SENTRYDISABLE;
    input CFGPOWERSTATECHANGEACK;
    input CFGREQPMTRANSITIONL23READY;
    input [7:0] CFGREVIDPF0;
    input [7:0] CFGREVIDPF1;
    input [7:0] CFGREVIDPF2;
    input [7:0] CFGREVIDPF3;
    input [15:0] CFGSUBSYSIDPF0;
    input [15:0] CFGSUBSYSIDPF1;
    input [15:0] CFGSUBSYSIDPF2;
    input [15:0] CFGSUBSYSIDPF3;
    input [15:0] CFGSUBSYSVENDID;
    input [35:0] CFGTPHRAMREADDATA;
    input [15:0] CFGVENDID;
    input CFGVFFLRDONE;
    input [7:0] CFGVFFLRFUNCNUM;
    input CONFMCAPREQUESTBYCONF;
    input [31:0] CONFREQDATA;
    input [3:0] CONFREQREGNUM;
    input [1:0] CONFREQTYPE;
    input CONFREQVALID;
    input CORECLK;
    input CORECLKCCIX;
    input CORECLKMIREPLAYRAM0;
    input CORECLKMIREPLAYRAM1;
    input CORECLKMIRXCOMPLETIONRAM0;
    input CORECLKMIRXCOMPLETIONRAM1;
    input CORECLKMIRXPOSTEDREQUESTRAM0;
    input CORECLKMIRXPOSTEDREQUESTRAM1;
    input [5:0] DBGSEL0;
    input [5:0] DBGSEL1;
    input [9:0] DRPADDR;
    input DRPCLK;
    input [15:0] DRPDI;
    input DRPEN;
    input DRPWE;
    input [21:0] MAXISCQTREADY;
    input [21:0] MAXISRCTREADY;
    input MCAPCLK;
    input MCAPPERST0B;
    input MCAPPERST1B;
    input MGMTRESETN;
    input MGMTSTICKYRESETN;
    input [5:0] MIREPLAYRAMERRCOR;
    input [5:0] MIREPLAYRAMERRUNCOR;
    input [127:0] MIREPLAYRAMREADDATA0;
    input [127:0] MIREPLAYRAMREADDATA1;
    input [11:0] MIRXCOMPLETIONRAMERRCOR;
    input [11:0] MIRXCOMPLETIONRAMERRUNCOR;
    input [143:0] MIRXCOMPLETIONRAMREADDATA0;
    input [143:0] MIRXCOMPLETIONRAMREADDATA1;
    input [5:0] MIRXPOSTEDREQUESTRAMERRCOR;
    input [5:0] MIRXPOSTEDREQUESTRAMERRUNCOR;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA0;
    input [143:0] MIRXPOSTEDREQUESTRAMREADDATA1;
    input [1:0] PCIECOMPLDELIVERED;
    input [7:0] PCIECOMPLDELIVEREDTAG0;
    input [7:0] PCIECOMPLDELIVEREDTAG1;
    input [1:0] PCIECQNPREQ;
    input PCIECQNPUSERCREDITRCVD;
    input PCIECQPIPELINEEMPTY;
    input PCIEPOSTEDREQDELIVERED;
    input PIPECLK;
    input PIPECLKEN;
    input [5:0] PIPEEQFS;
    input [5:0] PIPEEQLF;
    input PIPERESETN;
    input [1:0] PIPERX00CHARISK;
    input [31:0] PIPERX00DATA;
    input PIPERX00DATAVALID;
    input PIPERX00ELECIDLE;
    input PIPERX00EQDONE;
    input PIPERX00EQLPADAPTDONE;
    input PIPERX00EQLPLFFSSEL;
    input [17:0] PIPERX00EQLPNEWTXCOEFFORPRESET;
    input PIPERX00PHYSTATUS;
    input [1:0] PIPERX00STARTBLOCK;
    input [2:0] PIPERX00STATUS;
    input [1:0] PIPERX00SYNCHEADER;
    input PIPERX00VALID;
    input [1:0] PIPERX01CHARISK;
    input [31:0] PIPERX01DATA;
    input PIPERX01DATAVALID;
    input PIPERX01ELECIDLE;
    input PIPERX01EQDONE;
    input PIPERX01EQLPADAPTDONE;
    input PIPERX01EQLPLFFSSEL;
    input [17:0] PIPERX01EQLPNEWTXCOEFFORPRESET;
    input PIPERX01PHYSTATUS;
    input [1:0] PIPERX01STARTBLOCK;
    input [2:0] PIPERX01STATUS;
    input [1:0] PIPERX01SYNCHEADER;
    input PIPERX01VALID;
    input [1:0] PIPERX02CHARISK;
    input [31:0] PIPERX02DATA;
    input PIPERX02DATAVALID;
    input PIPERX02ELECIDLE;
    input PIPERX02EQDONE;
    input PIPERX02EQLPADAPTDONE;
    input PIPERX02EQLPLFFSSEL;
    input [17:0] PIPERX02EQLPNEWTXCOEFFORPRESET;
    input PIPERX02PHYSTATUS;
    input [1:0] PIPERX02STARTBLOCK;
    input [2:0] PIPERX02STATUS;
    input [1:0] PIPERX02SYNCHEADER;
    input PIPERX02VALID;
    input [1:0] PIPERX03CHARISK;
    input [31:0] PIPERX03DATA;
    input PIPERX03DATAVALID;
    input PIPERX03ELECIDLE;
    input PIPERX03EQDONE;
    input PIPERX03EQLPADAPTDONE;
    input PIPERX03EQLPLFFSSEL;
    input [17:0] PIPERX03EQLPNEWTXCOEFFORPRESET;
    input PIPERX03PHYSTATUS;
    input [1:0] PIPERX03STARTBLOCK;
    input [2:0] PIPERX03STATUS;
    input [1:0] PIPERX03SYNCHEADER;
    input PIPERX03VALID;
    input [1:0] PIPERX04CHARISK;
    input [31:0] PIPERX04DATA;
    input PIPERX04DATAVALID;
    input PIPERX04ELECIDLE;
    input PIPERX04EQDONE;
    input PIPERX04EQLPADAPTDONE;
    input PIPERX04EQLPLFFSSEL;
    input [17:0] PIPERX04EQLPNEWTXCOEFFORPRESET;
    input PIPERX04PHYSTATUS;
    input [1:0] PIPERX04STARTBLOCK;
    input [2:0] PIPERX04STATUS;
    input [1:0] PIPERX04SYNCHEADER;
    input PIPERX04VALID;
    input [1:0] PIPERX05CHARISK;
    input [31:0] PIPERX05DATA;
    input PIPERX05DATAVALID;
    input PIPERX05ELECIDLE;
    input PIPERX05EQDONE;
    input PIPERX05EQLPADAPTDONE;
    input PIPERX05EQLPLFFSSEL;
    input [17:0] PIPERX05EQLPNEWTXCOEFFORPRESET;
    input PIPERX05PHYSTATUS;
    input [1:0] PIPERX05STARTBLOCK;
    input [2:0] PIPERX05STATUS;
    input [1:0] PIPERX05SYNCHEADER;
    input PIPERX05VALID;
    input [1:0] PIPERX06CHARISK;
    input [31:0] PIPERX06DATA;
    input PIPERX06DATAVALID;
    input PIPERX06ELECIDLE;
    input PIPERX06EQDONE;
    input PIPERX06EQLPADAPTDONE;
    input PIPERX06EQLPLFFSSEL;
    input [17:0] PIPERX06EQLPNEWTXCOEFFORPRESET;
    input PIPERX06PHYSTATUS;
    input [1:0] PIPERX06STARTBLOCK;
    input [2:0] PIPERX06STATUS;
    input [1:0] PIPERX06SYNCHEADER;
    input PIPERX06VALID;
    input [1:0] PIPERX07CHARISK;
    input [31:0] PIPERX07DATA;
    input PIPERX07DATAVALID;
    input PIPERX07ELECIDLE;
    input PIPERX07EQDONE;
    input PIPERX07EQLPADAPTDONE;
    input PIPERX07EQLPLFFSSEL;
    input [17:0] PIPERX07EQLPNEWTXCOEFFORPRESET;
    input PIPERX07PHYSTATUS;
    input [1:0] PIPERX07STARTBLOCK;
    input [2:0] PIPERX07STATUS;
    input [1:0] PIPERX07SYNCHEADER;
    input PIPERX07VALID;
    input [1:0] PIPERX08CHARISK;
    input [31:0] PIPERX08DATA;
    input PIPERX08DATAVALID;
    input PIPERX08ELECIDLE;
    input PIPERX08EQDONE;
    input PIPERX08EQLPADAPTDONE;
    input PIPERX08EQLPLFFSSEL;
    input [17:0] PIPERX08EQLPNEWTXCOEFFORPRESET;
    input PIPERX08PHYSTATUS;
    input [1:0] PIPERX08STARTBLOCK;
    input [2:0] PIPERX08STATUS;
    input [1:0] PIPERX08SYNCHEADER;
    input PIPERX08VALID;
    input [1:0] PIPERX09CHARISK;
    input [31:0] PIPERX09DATA;
    input PIPERX09DATAVALID;
    input PIPERX09ELECIDLE;
    input PIPERX09EQDONE;
    input PIPERX09EQLPADAPTDONE;
    input PIPERX09EQLPLFFSSEL;
    input [17:0] PIPERX09EQLPNEWTXCOEFFORPRESET;
    input PIPERX09PHYSTATUS;
    input [1:0] PIPERX09STARTBLOCK;
    input [2:0] PIPERX09STATUS;
    input [1:0] PIPERX09SYNCHEADER;
    input PIPERX09VALID;
    input [1:0] PIPERX10CHARISK;
    input [31:0] PIPERX10DATA;
    input PIPERX10DATAVALID;
    input PIPERX10ELECIDLE;
    input PIPERX10EQDONE;
    input PIPERX10EQLPADAPTDONE;
    input PIPERX10EQLPLFFSSEL;
    input [17:0] PIPERX10EQLPNEWTXCOEFFORPRESET;
    input PIPERX10PHYSTATUS;
    input [1:0] PIPERX10STARTBLOCK;
    input [2:0] PIPERX10STATUS;
    input [1:0] PIPERX10SYNCHEADER;
    input PIPERX10VALID;
    input [1:0] PIPERX11CHARISK;
    input [31:0] PIPERX11DATA;
    input PIPERX11DATAVALID;
    input PIPERX11ELECIDLE;
    input PIPERX11EQDONE;
    input PIPERX11EQLPADAPTDONE;
    input PIPERX11EQLPLFFSSEL;
    input [17:0] PIPERX11EQLPNEWTXCOEFFORPRESET;
    input PIPERX11PHYSTATUS;
    input [1:0] PIPERX11STARTBLOCK;
    input [2:0] PIPERX11STATUS;
    input [1:0] PIPERX11SYNCHEADER;
    input PIPERX11VALID;
    input [1:0] PIPERX12CHARISK;
    input [31:0] PIPERX12DATA;
    input PIPERX12DATAVALID;
    input PIPERX12ELECIDLE;
    input PIPERX12EQDONE;
    input PIPERX12EQLPADAPTDONE;
    input PIPERX12EQLPLFFSSEL;
    input [17:0] PIPERX12EQLPNEWTXCOEFFORPRESET;
    input PIPERX12PHYSTATUS;
    input [1:0] PIPERX12STARTBLOCK;
    input [2:0] PIPERX12STATUS;
    input [1:0] PIPERX12SYNCHEADER;
    input PIPERX12VALID;
    input [1:0] PIPERX13CHARISK;
    input [31:0] PIPERX13DATA;
    input PIPERX13DATAVALID;
    input PIPERX13ELECIDLE;
    input PIPERX13EQDONE;
    input PIPERX13EQLPADAPTDONE;
    input PIPERX13EQLPLFFSSEL;
    input [17:0] PIPERX13EQLPNEWTXCOEFFORPRESET;
    input PIPERX13PHYSTATUS;
    input [1:0] PIPERX13STARTBLOCK;
    input [2:0] PIPERX13STATUS;
    input [1:0] PIPERX13SYNCHEADER;
    input PIPERX13VALID;
    input [1:0] PIPERX14CHARISK;
    input [31:0] PIPERX14DATA;
    input PIPERX14DATAVALID;
    input PIPERX14ELECIDLE;
    input PIPERX14EQDONE;
    input PIPERX14EQLPADAPTDONE;
    input PIPERX14EQLPLFFSSEL;
    input [17:0] PIPERX14EQLPNEWTXCOEFFORPRESET;
    input PIPERX14PHYSTATUS;
    input [1:0] PIPERX14STARTBLOCK;
    input [2:0] PIPERX14STATUS;
    input [1:0] PIPERX14SYNCHEADER;
    input PIPERX14VALID;
    input [1:0] PIPERX15CHARISK;
    input [31:0] PIPERX15DATA;
    input PIPERX15DATAVALID;
    input PIPERX15ELECIDLE;
    input PIPERX15EQDONE;
    input PIPERX15EQLPADAPTDONE;
    input PIPERX15EQLPLFFSSEL;
    input [17:0] PIPERX15EQLPNEWTXCOEFFORPRESET;
    input PIPERX15PHYSTATUS;
    input [1:0] PIPERX15STARTBLOCK;
    input [2:0] PIPERX15STATUS;
    input [1:0] PIPERX15SYNCHEADER;
    input PIPERX15VALID;
    input [17:0] PIPETX00EQCOEFF;
    input PIPETX00EQDONE;
    input [17:0] PIPETX01EQCOEFF;
    input PIPETX01EQDONE;
    input [17:0] PIPETX02EQCOEFF;
    input PIPETX02EQDONE;
    input [17:0] PIPETX03EQCOEFF;
    input PIPETX03EQDONE;
    input [17:0] PIPETX04EQCOEFF;
    input PIPETX04EQDONE;
    input [17:0] PIPETX05EQCOEFF;
    input PIPETX05EQDONE;
    input [17:0] PIPETX06EQCOEFF;
    input PIPETX06EQDONE;
    input [17:0] PIPETX07EQCOEFF;
    input PIPETX07EQDONE;
    input [17:0] PIPETX08EQCOEFF;
    input PIPETX08EQDONE;
    input [17:0] PIPETX09EQCOEFF;
    input PIPETX09EQDONE;
    input [17:0] PIPETX10EQCOEFF;
    input PIPETX10EQDONE;
    input [17:0] PIPETX11EQCOEFF;
    input PIPETX11EQDONE;
    input [17:0] PIPETX12EQCOEFF;
    input PIPETX12EQDONE;
    input [17:0] PIPETX13EQCOEFF;
    input PIPETX13EQDONE;
    input [17:0] PIPETX14EQCOEFF;
    input PIPETX14EQDONE;
    input [17:0] PIPETX15EQCOEFF;
    input PIPETX15EQDONE;
    input PLEQRESETEIEOSCOUNT;
    input PLGEN2UPSTREAMPREFERDEEMPH;
    input PLGEN34REDOEQSPEED;
    input PLGEN34REDOEQUALIZATION;
    input RESETN;
    input [255:0] SAXISCCIXTXTDATA;
    input [45:0] SAXISCCIXTXTUSER;
    input SAXISCCIXTXTVALID;
    input [255:0] SAXISCCTDATA;
    input [7:0] SAXISCCTKEEP;
    input SAXISCCTLAST;
    input [32:0] SAXISCCTUSER;
    input SAXISCCTVALID;
    input [255:0] SAXISRQTDATA;
    input [7:0] SAXISRQTKEEP;
    input SAXISRQTLAST;
    input [61:0] SAXISRQTUSER;
    input SAXISRQTVALID;
    input USERCLK;
    input USERCLK2;
    input USERCLKEN;
    input [31:0] USERSPAREIN;
endmodule

module TEMAC_SINGLE (...);
    parameter EMAC_1000BASEX_ENABLE = "FALSE";
    parameter EMAC_ADDRFILTER_ENABLE = "FALSE";
    parameter EMAC_BYTEPHY = "FALSE";
    parameter EMAC_CTRLLENCHECK_DISABLE = "FALSE";
    parameter [0:7] EMAC_DCRBASEADDR = 8'h00;
    parameter EMAC_GTLOOPBACK = "FALSE";
    parameter EMAC_HOST_ENABLE = "FALSE";
    parameter [8:0] EMAC_LINKTIMERVAL = 9'h000;
    parameter EMAC_LTCHECK_DISABLE = "FALSE";
    parameter EMAC_MDIO_ENABLE = "FALSE";
    parameter EMAC_MDIO_IGNORE_PHYADZERO = "FALSE";
    parameter [47:0] EMAC_PAUSEADDR = 48'h000000000000;
    parameter EMAC_PHYINITAUTONEG_ENABLE = "FALSE";
    parameter EMAC_PHYISOLATE = "FALSE";
    parameter EMAC_PHYLOOPBACKMSB = "FALSE";
    parameter EMAC_PHYPOWERDOWN = "FALSE";
    parameter EMAC_PHYRESET = "FALSE";
    parameter EMAC_RGMII_ENABLE = "FALSE";
    parameter EMAC_RX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_RXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_RXHALFDUPLEX = "FALSE";
    parameter EMAC_RXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_RXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_RXRESET = "FALSE";
    parameter EMAC_RXVLAN_ENABLE = "FALSE";
    parameter EMAC_RX_ENABLE = "TRUE";
    parameter EMAC_SGMII_ENABLE = "FALSE";
    parameter EMAC_SPEED_LSB = "FALSE";
    parameter EMAC_SPEED_MSB = "FALSE";
    parameter EMAC_TX16BITCLIENT_ENABLE = "FALSE";
    parameter EMAC_TXFLOWCTRL_ENABLE = "FALSE";
    parameter EMAC_TXHALFDUPLEX = "FALSE";
    parameter EMAC_TXIFGADJUST_ENABLE = "FALSE";
    parameter EMAC_TXINBANDFCS_ENABLE = "FALSE";
    parameter EMAC_TXJUMBOFRAME_ENABLE = "FALSE";
    parameter EMAC_TXRESET = "FALSE";
    parameter EMAC_TXVLAN_ENABLE = "FALSE";
    parameter EMAC_TX_ENABLE = "TRUE";
    parameter [47:0] EMAC_UNICASTADDR = 48'h000000000000;
    parameter EMAC_UNIDIRECTION_ENABLE = "FALSE";
    parameter EMAC_USECLKEN = "FALSE";
    parameter SIM_VERSION = "1.0";
    output DCRHOSTDONEIR;
    output EMACCLIENTANINTERRUPT;
    output EMACCLIENTRXBADFRAME;
    output EMACCLIENTRXCLIENTCLKOUT;
    output EMACCLIENTRXDVLD;
    output EMACCLIENTRXDVLDMSW;
    output EMACCLIENTRXFRAMEDROP;
    output EMACCLIENTRXGOODFRAME;
    output EMACCLIENTRXSTATSBYTEVLD;
    output EMACCLIENTRXSTATSVLD;
    output EMACCLIENTTXACK;
    output EMACCLIENTTXCLIENTCLKOUT;
    output EMACCLIENTTXCOLLISION;
    output EMACCLIENTTXRETRANSMIT;
    output EMACCLIENTTXSTATS;
    output EMACCLIENTTXSTATSBYTEVLD;
    output EMACCLIENTTXSTATSVLD;
    output EMACDCRACK;
    output EMACPHYENCOMMAALIGN;
    output EMACPHYLOOPBACKMSB;
    output EMACPHYMCLKOUT;
    output EMACPHYMDOUT;
    output EMACPHYMDTRI;
    output EMACPHYMGTRXRESET;
    output EMACPHYMGTTXRESET;
    output EMACPHYPOWERDOWN;
    output EMACPHYSYNCACQSTATUS;
    output EMACPHYTXCHARDISPMODE;
    output EMACPHYTXCHARDISPVAL;
    output EMACPHYTXCHARISK;
    output EMACPHYTXCLK;
    output EMACPHYTXEN;
    output EMACPHYTXER;
    output EMACPHYTXGMIIMIICLKOUT;
    output EMACSPEEDIS10100;
    output HOSTMIIMRDY;
    output [0:31] EMACDCRDBUS;
    output [15:0] EMACCLIENTRXD;
    output [31:0] HOSTRDDATA;
    output [6:0] EMACCLIENTRXSTATS;
    output [7:0] EMACPHYTXD;
    input CLIENTEMACDCMLOCKED;
    input CLIENTEMACPAUSEREQ;
    input CLIENTEMACRXCLIENTCLKIN;
    input CLIENTEMACTXCLIENTCLKIN;
    input CLIENTEMACTXDVLD;
    input CLIENTEMACTXDVLDMSW;
    input CLIENTEMACTXFIRSTBYTE;
    input CLIENTEMACTXUNDERRUN;
    input DCREMACCLK;
    input DCREMACENABLE;
    input DCREMACREAD;
    input DCREMACWRITE;
    input HOSTCLK;
    input HOSTMIIMSEL;
    input HOSTREQ;
    input PHYEMACCOL;
    input PHYEMACCRS;
    input PHYEMACGTXCLK;
    input PHYEMACMCLKIN;
    input PHYEMACMDIN;
    input PHYEMACMIITXCLK;
    input PHYEMACRXCHARISCOMMA;
    input PHYEMACRXCHARISK;
    input PHYEMACRXCLK;
    input PHYEMACRXDISPERR;
    input PHYEMACRXDV;
    input PHYEMACRXER;
    input PHYEMACRXNOTINTABLE;
    input PHYEMACRXRUNDISP;
    input PHYEMACSIGNALDET;
    input PHYEMACTXBUFERR;
    input PHYEMACTXGMIIMIICLKIN;
    input RESET;
    input [0:31] DCREMACDBUS;
    input [0:9] DCREMACABUS;
    input [15:0] CLIENTEMACPAUSEVAL;
    input [15:0] CLIENTEMACTXD;
    input [1:0] HOSTOPCODE;
    input [1:0] PHYEMACRXBUFSTATUS;
    input [2:0] PHYEMACRXCLKCORCNT;
    input [31:0] HOSTWRDATA;
    input [4:0] PHYEMACPHYAD;
    input [7:0] CLIENTEMACTXIFGDELAY;
    input [7:0] PHYEMACRXD;
    input [9:0] HOSTADDR;
endmodule

module CMAC (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [6:0] STAT_RX_BAD_CODE;
    output [3:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [3:0] STAT_RX_FRAGMENT;
    output [3:0] STAT_RX_FRAMING_ERR_0;
    output [3:0] STAT_RX_FRAMING_ERR_1;
    output [3:0] STAT_RX_FRAMING_ERR_10;
    output [3:0] STAT_RX_FRAMING_ERR_11;
    output [3:0] STAT_RX_FRAMING_ERR_12;
    output [3:0] STAT_RX_FRAMING_ERR_13;
    output [3:0] STAT_RX_FRAMING_ERR_14;
    output [3:0] STAT_RX_FRAMING_ERR_15;
    output [3:0] STAT_RX_FRAMING_ERR_16;
    output [3:0] STAT_RX_FRAMING_ERR_17;
    output [3:0] STAT_RX_FRAMING_ERR_18;
    output [3:0] STAT_RX_FRAMING_ERR_19;
    output [3:0] STAT_RX_FRAMING_ERR_2;
    output [3:0] STAT_RX_FRAMING_ERR_3;
    output [3:0] STAT_RX_FRAMING_ERR_4;
    output [3:0] STAT_RX_FRAMING_ERR_5;
    output [3:0] STAT_RX_FRAMING_ERR_6;
    output [3:0] STAT_RX_FRAMING_ERR_7;
    output [3:0] STAT_RX_FRAMING_ERR_8;
    output [3:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [3:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_STATUS;
    output [3:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [7:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [3:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [3:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [6:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module CMACE4 (...);
    parameter CTL_PTP_TRANSPCLK_MODE = "FALSE";
    parameter CTL_RX_CHECK_ACK = "TRUE";
    parameter CTL_RX_CHECK_PREAMBLE = "FALSE";
    parameter CTL_RX_CHECK_SFD = "FALSE";
    parameter CTL_RX_DELETE_FCS = "TRUE";
    parameter [15:0] CTL_RX_ETYPE_GCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_GPP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PCP = 16'h8808;
    parameter [15:0] CTL_RX_ETYPE_PPP = 16'h8808;
    parameter CTL_RX_FORWARD_CONTROL = "FALSE";
    parameter CTL_RX_IGNORE_FCS = "FALSE";
    parameter [14:0] CTL_RX_MAX_PACKET_LEN = 15'h2580;
    parameter [7:0] CTL_RX_MIN_PACKET_LEN = 8'h40;
    parameter [15:0] CTL_RX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_RX_OPCODE_MAX_GCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MAX_PCP = 16'hFFFF;
    parameter [15:0] CTL_RX_OPCODE_MIN_GCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_MIN_PCP = 16'h0000;
    parameter [15:0] CTL_RX_OPCODE_PPP = 16'h0001;
    parameter [47:0] CTL_RX_PAUSE_DA_MCAST = 48'h0180C2000001;
    parameter [47:0] CTL_RX_PAUSE_DA_UCAST = 48'h000000000000;
    parameter [47:0] CTL_RX_PAUSE_SA = 48'h000000000000;
    parameter CTL_RX_PROCESS_LFI = "FALSE";
    parameter [8:0] CTL_RX_RSFEC_AM_THRESHOLD = 9'h046;
    parameter [1:0] CTL_RX_RSFEC_FILL_ADJUST = 2'h0;
    parameter [15:0] CTL_RX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_RX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_RX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_RX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_RX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_RX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_RX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_RX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_RX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_RX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_RX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_RX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_RX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_RX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_RX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_RX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_RX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_RX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_RX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_RX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter CTL_TX_CUSTOM_PREAMBLE_ENABLE = "FALSE";
    parameter [47:0] CTL_TX_DA_GPP = 48'h0180C2000001;
    parameter [47:0] CTL_TX_DA_PPP = 48'h0180C2000001;
    parameter [15:0] CTL_TX_ETHERTYPE_GPP = 16'h8808;
    parameter [15:0] CTL_TX_ETHERTYPE_PPP = 16'h8808;
    parameter CTL_TX_FCS_INS_ENABLE = "TRUE";
    parameter CTL_TX_IGNORE_FCS = "FALSE";
    parameter [3:0] CTL_TX_IPG_VALUE = 4'hC;
    parameter [15:0] CTL_TX_OPCODE_GPP = 16'h0001;
    parameter [15:0] CTL_TX_OPCODE_PPP = 16'h0001;
    parameter CTL_TX_PTP_1STEP_ENABLE = "FALSE";
    parameter [10:0] CTL_TX_PTP_LATENCY_ADJUST = 11'h2C1;
    parameter [47:0] CTL_TX_SA_GPP = 48'h000000000000;
    parameter [47:0] CTL_TX_SA_PPP = 48'h000000000000;
    parameter [15:0] CTL_TX_VL_LENGTH_MINUS1 = 16'h3FFF;
    parameter [63:0] CTL_TX_VL_MARKER_ID0 = 64'hC16821003E97DE00;
    parameter [63:0] CTL_TX_VL_MARKER_ID1 = 64'h9D718E00628E7100;
    parameter [63:0] CTL_TX_VL_MARKER_ID10 = 64'hFD6C990002936600;
    parameter [63:0] CTL_TX_VL_MARKER_ID11 = 64'hB9915500466EAA00;
    parameter [63:0] CTL_TX_VL_MARKER_ID12 = 64'h5CB9B200A3464D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID13 = 64'h1AF8BD00E5074200;
    parameter [63:0] CTL_TX_VL_MARKER_ID14 = 64'h83C7CA007C383500;
    parameter [63:0] CTL_TX_VL_MARKER_ID15 = 64'h3536CD00CAC93200;
    parameter [63:0] CTL_TX_VL_MARKER_ID16 = 64'hC4314C003BCEB300;
    parameter [63:0] CTL_TX_VL_MARKER_ID17 = 64'hADD6B70052294800;
    parameter [63:0] CTL_TX_VL_MARKER_ID18 = 64'h5F662A00A099D500;
    parameter [63:0] CTL_TX_VL_MARKER_ID19 = 64'hC0F0E5003F0F1A00;
    parameter [63:0] CTL_TX_VL_MARKER_ID2 = 64'h594BE800A6B41700;
    parameter [63:0] CTL_TX_VL_MARKER_ID3 = 64'h4D957B00B26A8400;
    parameter [63:0] CTL_TX_VL_MARKER_ID4 = 64'hF50709000AF8F600;
    parameter [63:0] CTL_TX_VL_MARKER_ID5 = 64'hDD14C20022EB3D00;
    parameter [63:0] CTL_TX_VL_MARKER_ID6 = 64'h9A4A260065B5D900;
    parameter [63:0] CTL_TX_VL_MARKER_ID7 = 64'h7B45660084BA9900;
    parameter [63:0] CTL_TX_VL_MARKER_ID8 = 64'hA02476005FDB8900;
    parameter [63:0] CTL_TX_VL_MARKER_ID9 = 64'h68C9FB0097360400;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [329:0] RSFEC_BYPASS_RX_DOUT;
    output RSFEC_BYPASS_RX_DOUT_CW_START;
    output RSFEC_BYPASS_RX_DOUT_VALID;
    output [329:0] RSFEC_BYPASS_TX_DOUT;
    output RSFEC_BYPASS_TX_DOUT_CW_START;
    output RSFEC_BYPASS_TX_DOUT_VALID;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [6:0] RX_LANE_ALIGNER_FILL_0;
    output [6:0] RX_LANE_ALIGNER_FILL_1;
    output [6:0] RX_LANE_ALIGNER_FILL_10;
    output [6:0] RX_LANE_ALIGNER_FILL_11;
    output [6:0] RX_LANE_ALIGNER_FILL_12;
    output [6:0] RX_LANE_ALIGNER_FILL_13;
    output [6:0] RX_LANE_ALIGNER_FILL_14;
    output [6:0] RX_LANE_ALIGNER_FILL_15;
    output [6:0] RX_LANE_ALIGNER_FILL_16;
    output [6:0] RX_LANE_ALIGNER_FILL_17;
    output [6:0] RX_LANE_ALIGNER_FILL_18;
    output [6:0] RX_LANE_ALIGNER_FILL_19;
    output [6:0] RX_LANE_ALIGNER_FILL_2;
    output [6:0] RX_LANE_ALIGNER_FILL_3;
    output [6:0] RX_LANE_ALIGNER_FILL_4;
    output [6:0] RX_LANE_ALIGNER_FILL_5;
    output [6:0] RX_LANE_ALIGNER_FILL_6;
    output [6:0] RX_LANE_ALIGNER_FILL_7;
    output [6:0] RX_LANE_ALIGNER_FILL_8;
    output [6:0] RX_LANE_ALIGNER_FILL_9;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output [7:0] RX_OTN_BIP8_0;
    output [7:0] RX_OTN_BIP8_1;
    output [7:0] RX_OTN_BIP8_2;
    output [7:0] RX_OTN_BIP8_3;
    output [7:0] RX_OTN_BIP8_4;
    output [65:0] RX_OTN_DATA_0;
    output [65:0] RX_OTN_DATA_1;
    output [65:0] RX_OTN_DATA_2;
    output [65:0] RX_OTN_DATA_3;
    output [65:0] RX_OTN_DATA_4;
    output RX_OTN_ENA;
    output RX_OTN_LANE0;
    output RX_OTN_VLMARKER;
    output [55:0] RX_PREOUT;
    output [4:0] RX_PTP_PCSLANE_OUT;
    output [79:0] RX_PTP_TSTAMP_OUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [2:0] STAT_RX_BAD_CODE;
    output [2:0] STAT_RX_BAD_FCS;
    output STAT_RX_BAD_PREAMBLE;
    output STAT_RX_BAD_SFD;
    output STAT_RX_BIP_ERR_0;
    output STAT_RX_BIP_ERR_1;
    output STAT_RX_BIP_ERR_10;
    output STAT_RX_BIP_ERR_11;
    output STAT_RX_BIP_ERR_12;
    output STAT_RX_BIP_ERR_13;
    output STAT_RX_BIP_ERR_14;
    output STAT_RX_BIP_ERR_15;
    output STAT_RX_BIP_ERR_16;
    output STAT_RX_BIP_ERR_17;
    output STAT_RX_BIP_ERR_18;
    output STAT_RX_BIP_ERR_19;
    output STAT_RX_BIP_ERR_2;
    output STAT_RX_BIP_ERR_3;
    output STAT_RX_BIP_ERR_4;
    output STAT_RX_BIP_ERR_5;
    output STAT_RX_BIP_ERR_6;
    output STAT_RX_BIP_ERR_7;
    output STAT_RX_BIP_ERR_8;
    output STAT_RX_BIP_ERR_9;
    output [19:0] STAT_RX_BLOCK_LOCK;
    output STAT_RX_BROADCAST;
    output [2:0] STAT_RX_FRAGMENT;
    output [1:0] STAT_RX_FRAMING_ERR_0;
    output [1:0] STAT_RX_FRAMING_ERR_1;
    output [1:0] STAT_RX_FRAMING_ERR_10;
    output [1:0] STAT_RX_FRAMING_ERR_11;
    output [1:0] STAT_RX_FRAMING_ERR_12;
    output [1:0] STAT_RX_FRAMING_ERR_13;
    output [1:0] STAT_RX_FRAMING_ERR_14;
    output [1:0] STAT_RX_FRAMING_ERR_15;
    output [1:0] STAT_RX_FRAMING_ERR_16;
    output [1:0] STAT_RX_FRAMING_ERR_17;
    output [1:0] STAT_RX_FRAMING_ERR_18;
    output [1:0] STAT_RX_FRAMING_ERR_19;
    output [1:0] STAT_RX_FRAMING_ERR_2;
    output [1:0] STAT_RX_FRAMING_ERR_3;
    output [1:0] STAT_RX_FRAMING_ERR_4;
    output [1:0] STAT_RX_FRAMING_ERR_5;
    output [1:0] STAT_RX_FRAMING_ERR_6;
    output [1:0] STAT_RX_FRAMING_ERR_7;
    output [1:0] STAT_RX_FRAMING_ERR_8;
    output [1:0] STAT_RX_FRAMING_ERR_9;
    output STAT_RX_FRAMING_ERR_VALID_0;
    output STAT_RX_FRAMING_ERR_VALID_1;
    output STAT_RX_FRAMING_ERR_VALID_10;
    output STAT_RX_FRAMING_ERR_VALID_11;
    output STAT_RX_FRAMING_ERR_VALID_12;
    output STAT_RX_FRAMING_ERR_VALID_13;
    output STAT_RX_FRAMING_ERR_VALID_14;
    output STAT_RX_FRAMING_ERR_VALID_15;
    output STAT_RX_FRAMING_ERR_VALID_16;
    output STAT_RX_FRAMING_ERR_VALID_17;
    output STAT_RX_FRAMING_ERR_VALID_18;
    output STAT_RX_FRAMING_ERR_VALID_19;
    output STAT_RX_FRAMING_ERR_VALID_2;
    output STAT_RX_FRAMING_ERR_VALID_3;
    output STAT_RX_FRAMING_ERR_VALID_4;
    output STAT_RX_FRAMING_ERR_VALID_5;
    output STAT_RX_FRAMING_ERR_VALID_6;
    output STAT_RX_FRAMING_ERR_VALID_7;
    output STAT_RX_FRAMING_ERR_VALID_8;
    output STAT_RX_FRAMING_ERR_VALID_9;
    output STAT_RX_GOT_SIGNAL_OS;
    output STAT_RX_HI_BER;
    output STAT_RX_INRANGEERR;
    output STAT_RX_INTERNAL_LOCAL_FAULT;
    output STAT_RX_JABBER;
    output [7:0] STAT_RX_LANE0_VLM_BIP7;
    output STAT_RX_LANE0_VLM_BIP7_VALID;
    output STAT_RX_LOCAL_FAULT;
    output [19:0] STAT_RX_MF_ERR;
    output [19:0] STAT_RX_MF_LEN_ERR;
    output [19:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MULTICAST;
    output STAT_RX_OVERSIZE;
    output STAT_RX_PACKET_1024_1518_BYTES;
    output STAT_RX_PACKET_128_255_BYTES;
    output STAT_RX_PACKET_1519_1522_BYTES;
    output STAT_RX_PACKET_1523_1548_BYTES;
    output STAT_RX_PACKET_1549_2047_BYTES;
    output STAT_RX_PACKET_2048_4095_BYTES;
    output STAT_RX_PACKET_256_511_BYTES;
    output STAT_RX_PACKET_4096_8191_BYTES;
    output STAT_RX_PACKET_512_1023_BYTES;
    output STAT_RX_PACKET_64_BYTES;
    output STAT_RX_PACKET_65_127_BYTES;
    output STAT_RX_PACKET_8192_9215_BYTES;
    output STAT_RX_PACKET_BAD_FCS;
    output STAT_RX_PACKET_LARGE;
    output [2:0] STAT_RX_PACKET_SMALL;
    output STAT_RX_PAUSE;
    output [15:0] STAT_RX_PAUSE_QUANTA0;
    output [15:0] STAT_RX_PAUSE_QUANTA1;
    output [15:0] STAT_RX_PAUSE_QUANTA2;
    output [15:0] STAT_RX_PAUSE_QUANTA3;
    output [15:0] STAT_RX_PAUSE_QUANTA4;
    output [15:0] STAT_RX_PAUSE_QUANTA5;
    output [15:0] STAT_RX_PAUSE_QUANTA6;
    output [15:0] STAT_RX_PAUSE_QUANTA7;
    output [15:0] STAT_RX_PAUSE_QUANTA8;
    output [8:0] STAT_RX_PAUSE_REQ;
    output [8:0] STAT_RX_PAUSE_VALID;
    output STAT_RX_RECEIVED_LOCAL_FAULT;
    output STAT_RX_REMOTE_FAULT;
    output STAT_RX_RSFEC_AM_LOCK0;
    output STAT_RX_RSFEC_AM_LOCK1;
    output STAT_RX_RSFEC_AM_LOCK2;
    output STAT_RX_RSFEC_AM_LOCK3;
    output STAT_RX_RSFEC_CORRECTED_CW_INC;
    output STAT_RX_RSFEC_CW_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT0_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT1_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT2_INC;
    output [2:0] STAT_RX_RSFEC_ERR_COUNT3_INC;
    output STAT_RX_RSFEC_HI_SER;
    output STAT_RX_RSFEC_LANE_ALIGNMENT_STATUS;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_0;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_1;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_2;
    output [13:0] STAT_RX_RSFEC_LANE_FILL_3;
    output [7:0] STAT_RX_RSFEC_LANE_MAPPING;
    output [31:0] STAT_RX_RSFEC_RSVD;
    output STAT_RX_RSFEC_UNCORRECTED_CW_INC;
    output STAT_RX_STATUS;
    output [2:0] STAT_RX_STOMPED_FCS;
    output [19:0] STAT_RX_SYNCED;
    output [19:0] STAT_RX_SYNCED_ERR;
    output [2:0] STAT_RX_TEST_PATTERN_MISMATCH;
    output STAT_RX_TOOLONG;
    output [6:0] STAT_RX_TOTAL_BYTES;
    output [13:0] STAT_RX_TOTAL_GOOD_BYTES;
    output STAT_RX_TOTAL_GOOD_PACKETS;
    output [2:0] STAT_RX_TOTAL_PACKETS;
    output STAT_RX_TRUNCATED;
    output [2:0] STAT_RX_UNDERSIZE;
    output STAT_RX_UNICAST;
    output STAT_RX_USER_PAUSE;
    output STAT_RX_VLAN;
    output [19:0] STAT_RX_VL_DEMUXED;
    output [4:0] STAT_RX_VL_NUMBER_0;
    output [4:0] STAT_RX_VL_NUMBER_1;
    output [4:0] STAT_RX_VL_NUMBER_10;
    output [4:0] STAT_RX_VL_NUMBER_11;
    output [4:0] STAT_RX_VL_NUMBER_12;
    output [4:0] STAT_RX_VL_NUMBER_13;
    output [4:0] STAT_RX_VL_NUMBER_14;
    output [4:0] STAT_RX_VL_NUMBER_15;
    output [4:0] STAT_RX_VL_NUMBER_16;
    output [4:0] STAT_RX_VL_NUMBER_17;
    output [4:0] STAT_RX_VL_NUMBER_18;
    output [4:0] STAT_RX_VL_NUMBER_19;
    output [4:0] STAT_RX_VL_NUMBER_2;
    output [4:0] STAT_RX_VL_NUMBER_3;
    output [4:0] STAT_RX_VL_NUMBER_4;
    output [4:0] STAT_RX_VL_NUMBER_5;
    output [4:0] STAT_RX_VL_NUMBER_6;
    output [4:0] STAT_RX_VL_NUMBER_7;
    output [4:0] STAT_RX_VL_NUMBER_8;
    output [4:0] STAT_RX_VL_NUMBER_9;
    output STAT_TX_BAD_FCS;
    output STAT_TX_BROADCAST;
    output STAT_TX_FRAME_ERROR;
    output STAT_TX_LOCAL_FAULT;
    output STAT_TX_MULTICAST;
    output STAT_TX_PACKET_1024_1518_BYTES;
    output STAT_TX_PACKET_128_255_BYTES;
    output STAT_TX_PACKET_1519_1522_BYTES;
    output STAT_TX_PACKET_1523_1548_BYTES;
    output STAT_TX_PACKET_1549_2047_BYTES;
    output STAT_TX_PACKET_2048_4095_BYTES;
    output STAT_TX_PACKET_256_511_BYTES;
    output STAT_TX_PACKET_4096_8191_BYTES;
    output STAT_TX_PACKET_512_1023_BYTES;
    output STAT_TX_PACKET_64_BYTES;
    output STAT_TX_PACKET_65_127_BYTES;
    output STAT_TX_PACKET_8192_9215_BYTES;
    output STAT_TX_PACKET_LARGE;
    output STAT_TX_PACKET_SMALL;
    output STAT_TX_PAUSE;
    output [8:0] STAT_TX_PAUSE_VALID;
    output STAT_TX_PTP_FIFO_READ_ERROR;
    output STAT_TX_PTP_FIFO_WRITE_ERROR;
    output [5:0] STAT_TX_TOTAL_BYTES;
    output [13:0] STAT_TX_TOTAL_GOOD_BYTES;
    output STAT_TX_TOTAL_GOOD_PACKETS;
    output STAT_TX_TOTAL_PACKETS;
    output STAT_TX_UNICAST;
    output STAT_TX_USER_PAUSE;
    output STAT_TX_VLAN;
    output TX_OVFOUT;
    output [4:0] TX_PTP_PCSLANE_OUT;
    output [79:0] TX_PTP_TSTAMP_OUT;
    output [15:0] TX_PTP_TSTAMP_TAG_OUT;
    output TX_PTP_TSTAMP_VALID_OUT;
    output TX_RDYOUT;
    output [15:0] TX_SERDES_ALT_DATA0;
    output [15:0] TX_SERDES_ALT_DATA1;
    output [15:0] TX_SERDES_ALT_DATA2;
    output [15:0] TX_SERDES_ALT_DATA3;
    output [63:0] TX_SERDES_DATA0;
    output [63:0] TX_SERDES_DATA1;
    output [63:0] TX_SERDES_DATA2;
    output [63:0] TX_SERDES_DATA3;
    output [31:0] TX_SERDES_DATA4;
    output [31:0] TX_SERDES_DATA5;
    output [31:0] TX_SERDES_DATA6;
    output [31:0] TX_SERDES_DATA7;
    output [31:0] TX_SERDES_DATA8;
    output [31:0] TX_SERDES_DATA9;
    output TX_UNFOUT;
    input CTL_CAUI4_MODE;
    input CTL_RSFEC_ENABLE_TRANSCODER_BYPASS_MODE;
    input CTL_RSFEC_IEEE_ERROR_INDICATION_MODE;
    input CTL_RX_CHECK_ETYPE_GCP;
    input CTL_RX_CHECK_ETYPE_GPP;
    input CTL_RX_CHECK_ETYPE_PCP;
    input CTL_RX_CHECK_ETYPE_PPP;
    input CTL_RX_CHECK_MCAST_GCP;
    input CTL_RX_CHECK_MCAST_GPP;
    input CTL_RX_CHECK_MCAST_PCP;
    input CTL_RX_CHECK_MCAST_PPP;
    input CTL_RX_CHECK_OPCODE_GCP;
    input CTL_RX_CHECK_OPCODE_GPP;
    input CTL_RX_CHECK_OPCODE_PCP;
    input CTL_RX_CHECK_OPCODE_PPP;
    input CTL_RX_CHECK_SA_GCP;
    input CTL_RX_CHECK_SA_GPP;
    input CTL_RX_CHECK_SA_PCP;
    input CTL_RX_CHECK_SA_PPP;
    input CTL_RX_CHECK_UCAST_GCP;
    input CTL_RX_CHECK_UCAST_GPP;
    input CTL_RX_CHECK_UCAST_PCP;
    input CTL_RX_CHECK_UCAST_PPP;
    input CTL_RX_ENABLE;
    input CTL_RX_ENABLE_GCP;
    input CTL_RX_ENABLE_GPP;
    input CTL_RX_ENABLE_PCP;
    input CTL_RX_ENABLE_PPP;
    input CTL_RX_FORCE_RESYNC;
    input [8:0] CTL_RX_PAUSE_ACK;
    input [8:0] CTL_RX_PAUSE_ENABLE;
    input CTL_RX_RSFEC_ENABLE;
    input CTL_RX_RSFEC_ENABLE_CORRECTION;
    input CTL_RX_RSFEC_ENABLE_INDICATION;
    input [79:0] CTL_RX_SYSTEMTIMERIN;
    input CTL_RX_TEST_PATTERN;
    input CTL_TX_ENABLE;
    input CTL_TX_LANE0_VLM_BIP7_OVERRIDE;
    input [7:0] CTL_TX_LANE0_VLM_BIP7_OVERRIDE_VALUE;
    input [8:0] CTL_TX_PAUSE_ENABLE;
    input [15:0] CTL_TX_PAUSE_QUANTA0;
    input [15:0] CTL_TX_PAUSE_QUANTA1;
    input [15:0] CTL_TX_PAUSE_QUANTA2;
    input [15:0] CTL_TX_PAUSE_QUANTA3;
    input [15:0] CTL_TX_PAUSE_QUANTA4;
    input [15:0] CTL_TX_PAUSE_QUANTA5;
    input [15:0] CTL_TX_PAUSE_QUANTA6;
    input [15:0] CTL_TX_PAUSE_QUANTA7;
    input [15:0] CTL_TX_PAUSE_QUANTA8;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER0;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER1;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER2;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER3;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER4;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER5;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER6;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER7;
    input [15:0] CTL_TX_PAUSE_REFRESH_TIMER8;
    input [8:0] CTL_TX_PAUSE_REQ;
    input CTL_TX_PTP_VLANE_ADJUST_MODE;
    input CTL_TX_RESEND_PAUSE;
    input CTL_TX_RSFEC_ENABLE;
    input CTL_TX_SEND_IDLE;
    input CTL_TX_SEND_LFI;
    input CTL_TX_SEND_RFI;
    input [79:0] CTL_TX_SYSTEMTIMERIN;
    input CTL_TX_TEST_PATTERN;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input [329:0] RSFEC_BYPASS_RX_DIN;
    input RSFEC_BYPASS_RX_DIN_CW_START;
    input [329:0] RSFEC_BYPASS_TX_DIN;
    input RSFEC_BYPASS_TX_DIN_CW_START;
    input RX_CLK;
    input RX_RESET;
    input [15:0] RX_SERDES_ALT_DATA0;
    input [15:0] RX_SERDES_ALT_DATA1;
    input [15:0] RX_SERDES_ALT_DATA2;
    input [15:0] RX_SERDES_ALT_DATA3;
    input [9:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA0;
    input [63:0] RX_SERDES_DATA1;
    input [63:0] RX_SERDES_DATA2;
    input [63:0] RX_SERDES_DATA3;
    input [31:0] RX_SERDES_DATA4;
    input [31:0] RX_SERDES_DATA5;
    input [31:0] RX_SERDES_DATA6;
    input [31:0] RX_SERDES_DATA7;
    input [31:0] RX_SERDES_DATA8;
    input [31:0] RX_SERDES_DATA9;
    input [9:0] RX_SERDES_RESET;
    input TX_CLK;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input [55:0] TX_PREIN;
    input [1:0] TX_PTP_1588OP_IN;
    input [15:0] TX_PTP_CHKSUM_OFFSET_IN;
    input [63:0] TX_PTP_RXTSTAMP_IN;
    input [15:0] TX_PTP_TAG_FIELD_IN;
    input [15:0] TX_PTP_TSTAMP_OFFSET_IN;
    input TX_PTP_UPD_CHKSUM_IN;
    input TX_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

(* keep *)
module HBM_REF_CLK (...);
    input REF_CLK;
endmodule

(* keep *)
module HBM_SNGLBLI_INTF_APB (...);
    parameter CLK_SEL = "FALSE";
    parameter [0:0] IS_PCLK_INVERTED = 1'b0;
    parameter [0:0] IS_PRESET_N_INVERTED = 1'b0;
    parameter MC_ENABLE = "FALSE";
    parameter PHY_ENABLE = "FALSE";
    parameter PHY_PCLK_INVERT = "FALSE";
    parameter SWITCH_ENABLE = "FALSE";
    output CATTRIP_PIPE;
    output [31:0] PRDATA_PIPE;
    output PREADY_PIPE;
    output PSLVERR_PIPE;
    output [2:0] TEMP_PIPE;
    input [21:0] PADDR;
    (* invertible_pin = "IS_PCLK_INVERTED" *)
    input PCLK;
    input PENABLE;
    (* invertible_pin = "IS_PRESET_N_INVERTED" *)
    input PRESET_N;
    input PSEL;
    input [31:0] PWDATA;
    input PWRITE;
endmodule

(* keep *)
module HBM_SNGLBLI_INTF_AXI (...);
    parameter CLK_SEL = "FALSE";
    parameter integer DATARATE = 1800;
    parameter [0:0] IS_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_ARESET_N_INVERTED = 1'b0;
    parameter MC_ENABLE = "FALSE";
    parameter integer PAGEHIT_PERCENT = 75;
    parameter PHY_ENABLE = "FALSE";
    parameter integer READ_PERCENT = 50;
    parameter SWITCH_ENABLE = "FALSE";
    parameter integer WRITE_PERCENT = 50;
    output ARREADY_PIPE;
    output AWREADY_PIPE;
    output [5:0] BID_PIPE;
    output [1:0] BRESP_PIPE;
    output BVALID_PIPE;
    output [1:0] DFI_AW_AERR_N_PIPE;
    output DFI_CLK_BUF;
    output DFI_CTRLUPD_ACK_PIPE;
    output [7:0] DFI_DBI_BYTE_DISABLE_PIPE;
    output [20:0] DFI_DW_RDDATA_DBI_PIPE;
    output [7:0] DFI_DW_RDDATA_DERR_PIPE;
    output [1:0] DFI_DW_RDDATA_PAR_VALID_PIPE;
    output [1:0] DFI_DW_RDDATA_VALID_PIPE;
    output DFI_INIT_COMPLETE_PIPE;
    output DFI_PHYUPD_REQ_PIPE;
    output DFI_PHYUPD_TYPE_PIPE;
    output DFI_PHY_LP_STATE_PIPE;
    output DFI_RST_N_BUF;
    output [5:0] MC_STATUS;
    output [7:0] PHY_STATUS;
    output [31:0] RDATA_PARITY_PIPE;
    output [255:0] RDATA_PIPE;
    output [5:0] RID_PIPE;
    output RLAST_PIPE;
    output [1:0] RRESP_PIPE;
    output RVALID_PIPE;
    output [5:0] STATUS;
    output WREADY_PIPE;
    (* invertible_pin = "IS_ACLK_INVERTED" *)
    input ACLK;
    input [36:0] ARADDR;
    input [1:0] ARBURST;
    (* invertible_pin = "IS_ARESET_N_INVERTED" *)
    input ARESET_N;
    input [5:0] ARID;
    input [3:0] ARLEN;
    input [2:0] ARSIZE;
    input ARVALID;
    input [36:0] AWADDR;
    input [1:0] AWBURST;
    input [5:0] AWID;
    input [3:0] AWLEN;
    input [2:0] AWSIZE;
    input AWVALID;
    input BREADY;
    input BSCAN_CK;
    input DFI_LP_PWR_X_REQ;
    input MBIST_EN;
    input RREADY;
    input [255:0] WDATA;
    input [31:0] WDATA_PARITY;
    input WLAST;
    input [31:0] WSTRB;
    input WVALID;
endmodule

(* keep *)
module HBM_ONE_STACK_INTF (...);
    parameter CLK_SEL_00 = "FALSE";
    parameter CLK_SEL_01 = "FALSE";
    parameter CLK_SEL_02 = "FALSE";
    parameter CLK_SEL_03 = "FALSE";
    parameter CLK_SEL_04 = "FALSE";
    parameter CLK_SEL_05 = "FALSE";
    parameter CLK_SEL_06 = "FALSE";
    parameter CLK_SEL_07 = "FALSE";
    parameter CLK_SEL_08 = "FALSE";
    parameter CLK_SEL_09 = "FALSE";
    parameter CLK_SEL_10 = "FALSE";
    parameter CLK_SEL_11 = "FALSE";
    parameter CLK_SEL_12 = "FALSE";
    parameter CLK_SEL_13 = "FALSE";
    parameter CLK_SEL_14 = "FALSE";
    parameter CLK_SEL_15 = "FALSE";
    parameter integer DATARATE_00 = 1800;
    parameter integer DATARATE_01 = 1800;
    parameter integer DATARATE_02 = 1800;
    parameter integer DATARATE_03 = 1800;
    parameter integer DATARATE_04 = 1800;
    parameter integer DATARATE_05 = 1800;
    parameter integer DATARATE_06 = 1800;
    parameter integer DATARATE_07 = 1800;
    parameter DA_LOCKOUT = "FALSE";
    parameter [0:0] IS_APB_0_PCLK_INVERTED = 1'b0;
    parameter [0:0] IS_APB_0_PRESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_00_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_00_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_01_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_01_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_02_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_02_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_03_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_03_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_04_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_04_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_05_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_05_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_06_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_06_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_07_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_07_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_08_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_08_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_09_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_09_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_10_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_10_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_11_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_11_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_12_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_12_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_13_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_13_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_14_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_14_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_15_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_15_ARESET_N_INVERTED = 1'b0;
    parameter MC_ENABLE_0 = "FALSE";
    parameter MC_ENABLE_1 = "FALSE";
    parameter MC_ENABLE_2 = "FALSE";
    parameter MC_ENABLE_3 = "FALSE";
    parameter MC_ENABLE_4 = "FALSE";
    parameter MC_ENABLE_5 = "FALSE";
    parameter MC_ENABLE_6 = "FALSE";
    parameter MC_ENABLE_7 = "FALSE";
    parameter MC_ENABLE_APB = "FALSE";
    parameter integer PAGEHIT_PERCENT_00 = 75;
    parameter PHY_ENABLE_00 = "FALSE";
    parameter PHY_ENABLE_01 = "FALSE";
    parameter PHY_ENABLE_02 = "FALSE";
    parameter PHY_ENABLE_03 = "FALSE";
    parameter PHY_ENABLE_04 = "FALSE";
    parameter PHY_ENABLE_05 = "FALSE";
    parameter PHY_ENABLE_06 = "FALSE";
    parameter PHY_ENABLE_07 = "FALSE";
    parameter PHY_ENABLE_08 = "FALSE";
    parameter PHY_ENABLE_09 = "FALSE";
    parameter PHY_ENABLE_10 = "FALSE";
    parameter PHY_ENABLE_11 = "FALSE";
    parameter PHY_ENABLE_12 = "FALSE";
    parameter PHY_ENABLE_13 = "FALSE";
    parameter PHY_ENABLE_14 = "FALSE";
    parameter PHY_ENABLE_15 = "FALSE";
    parameter PHY_ENABLE_APB = "FALSE";
    parameter PHY_PCLK_INVERT_01 = "FALSE";
    parameter integer READ_PERCENT_00 = 50;
    parameter integer READ_PERCENT_01 = 50;
    parameter integer READ_PERCENT_02 = 50;
    parameter integer READ_PERCENT_03 = 50;
    parameter integer READ_PERCENT_04 = 50;
    parameter integer READ_PERCENT_05 = 50;
    parameter integer READ_PERCENT_06 = 50;
    parameter integer READ_PERCENT_07 = 50;
    parameter integer READ_PERCENT_08 = 50;
    parameter integer READ_PERCENT_09 = 50;
    parameter integer READ_PERCENT_10 = 50;
    parameter integer READ_PERCENT_11 = 50;
    parameter integer READ_PERCENT_12 = 50;
    parameter integer READ_PERCENT_13 = 50;
    parameter integer READ_PERCENT_14 = 50;
    parameter integer READ_PERCENT_15 = 50;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter integer STACK_LOCATION = 0;
    parameter SWITCH_ENABLE = "FALSE";
    parameter integer WRITE_PERCENT_00 = 50;
    parameter integer WRITE_PERCENT_01 = 50;
    parameter integer WRITE_PERCENT_02 = 50;
    parameter integer WRITE_PERCENT_03 = 50;
    parameter integer WRITE_PERCENT_04 = 50;
    parameter integer WRITE_PERCENT_05 = 50;
    parameter integer WRITE_PERCENT_06 = 50;
    parameter integer WRITE_PERCENT_07 = 50;
    parameter integer WRITE_PERCENT_08 = 50;
    parameter integer WRITE_PERCENT_09 = 50;
    parameter integer WRITE_PERCENT_10 = 50;
    parameter integer WRITE_PERCENT_11 = 50;
    parameter integer WRITE_PERCENT_12 = 50;
    parameter integer WRITE_PERCENT_13 = 50;
    parameter integer WRITE_PERCENT_14 = 50;
    parameter integer WRITE_PERCENT_15 = 50;
    output [31:0] APB_0_PRDATA;
    output APB_0_PREADY;
    output APB_0_PSLVERR;
    output AXI_00_ARREADY;
    output AXI_00_AWREADY;
    output [5:0] AXI_00_BID;
    output [1:0] AXI_00_BRESP;
    output AXI_00_BVALID;
    output [1:0] AXI_00_DFI_AW_AERR_N;
    output AXI_00_DFI_CLK_BUF;
    output [7:0] AXI_00_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_00_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_00_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_00_DFI_DW_RDDATA_VALID;
    output AXI_00_DFI_INIT_COMPLETE;
    output AXI_00_DFI_PHYUPD_REQ;
    output AXI_00_DFI_PHY_LP_STATE;
    output AXI_00_DFI_RST_N_BUF;
    output [5:0] AXI_00_MC_STATUS;
    output [7:0] AXI_00_PHY_STATUS;
    output [255:0] AXI_00_RDATA;
    output [31:0] AXI_00_RDATA_PARITY;
    output [5:0] AXI_00_RID;
    output AXI_00_RLAST;
    output [1:0] AXI_00_RRESP;
    output AXI_00_RVALID;
    output AXI_00_WREADY;
    output AXI_01_ARREADY;
    output AXI_01_AWREADY;
    output [5:0] AXI_01_BID;
    output [1:0] AXI_01_BRESP;
    output AXI_01_BVALID;
    output [1:0] AXI_01_DFI_AW_AERR_N;
    output AXI_01_DFI_CLK_BUF;
    output [7:0] AXI_01_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_01_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_01_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_01_DFI_DW_RDDATA_VALID;
    output AXI_01_DFI_INIT_COMPLETE;
    output AXI_01_DFI_PHYUPD_REQ;
    output AXI_01_DFI_PHY_LP_STATE;
    output AXI_01_DFI_RST_N_BUF;
    output [255:0] AXI_01_RDATA;
    output [31:0] AXI_01_RDATA_PARITY;
    output [5:0] AXI_01_RID;
    output AXI_01_RLAST;
    output [1:0] AXI_01_RRESP;
    output AXI_01_RVALID;
    output AXI_01_WREADY;
    output AXI_02_ARREADY;
    output AXI_02_AWREADY;
    output [5:0] AXI_02_BID;
    output [1:0] AXI_02_BRESP;
    output AXI_02_BVALID;
    output [1:0] AXI_02_DFI_AW_AERR_N;
    output AXI_02_DFI_CLK_BUF;
    output [7:0] AXI_02_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_02_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_02_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_02_DFI_DW_RDDATA_VALID;
    output AXI_02_DFI_INIT_COMPLETE;
    output AXI_02_DFI_PHYUPD_REQ;
    output AXI_02_DFI_PHY_LP_STATE;
    output AXI_02_DFI_RST_N_BUF;
    output [5:0] AXI_02_MC_STATUS;
    output [7:0] AXI_02_PHY_STATUS;
    output [255:0] AXI_02_RDATA;
    output [31:0] AXI_02_RDATA_PARITY;
    output [5:0] AXI_02_RID;
    output AXI_02_RLAST;
    output [1:0] AXI_02_RRESP;
    output AXI_02_RVALID;
    output AXI_02_WREADY;
    output AXI_03_ARREADY;
    output AXI_03_AWREADY;
    output [5:0] AXI_03_BID;
    output [1:0] AXI_03_BRESP;
    output AXI_03_BVALID;
    output [1:0] AXI_03_DFI_AW_AERR_N;
    output AXI_03_DFI_CLK_BUF;
    output [7:0] AXI_03_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_03_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_03_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_03_DFI_DW_RDDATA_VALID;
    output AXI_03_DFI_INIT_COMPLETE;
    output AXI_03_DFI_PHYUPD_REQ;
    output AXI_03_DFI_PHY_LP_STATE;
    output AXI_03_DFI_RST_N_BUF;
    output [255:0] AXI_03_RDATA;
    output [31:0] AXI_03_RDATA_PARITY;
    output [5:0] AXI_03_RID;
    output AXI_03_RLAST;
    output [1:0] AXI_03_RRESP;
    output AXI_03_RVALID;
    output AXI_03_WREADY;
    output AXI_04_ARREADY;
    output AXI_04_AWREADY;
    output [5:0] AXI_04_BID;
    output [1:0] AXI_04_BRESP;
    output AXI_04_BVALID;
    output [1:0] AXI_04_DFI_AW_AERR_N;
    output AXI_04_DFI_CLK_BUF;
    output [7:0] AXI_04_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_04_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_04_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_04_DFI_DW_RDDATA_VALID;
    output AXI_04_DFI_INIT_COMPLETE;
    output AXI_04_DFI_PHYUPD_REQ;
    output AXI_04_DFI_PHY_LP_STATE;
    output AXI_04_DFI_RST_N_BUF;
    output [5:0] AXI_04_MC_STATUS;
    output [7:0] AXI_04_PHY_STATUS;
    output [255:0] AXI_04_RDATA;
    output [31:0] AXI_04_RDATA_PARITY;
    output [5:0] AXI_04_RID;
    output AXI_04_RLAST;
    output [1:0] AXI_04_RRESP;
    output AXI_04_RVALID;
    output AXI_04_WREADY;
    output AXI_05_ARREADY;
    output AXI_05_AWREADY;
    output [5:0] AXI_05_BID;
    output [1:0] AXI_05_BRESP;
    output AXI_05_BVALID;
    output [1:0] AXI_05_DFI_AW_AERR_N;
    output AXI_05_DFI_CLK_BUF;
    output [7:0] AXI_05_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_05_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_05_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_05_DFI_DW_RDDATA_VALID;
    output AXI_05_DFI_INIT_COMPLETE;
    output AXI_05_DFI_PHYUPD_REQ;
    output AXI_05_DFI_PHY_LP_STATE;
    output AXI_05_DFI_RST_N_BUF;
    output [255:0] AXI_05_RDATA;
    output [31:0] AXI_05_RDATA_PARITY;
    output [5:0] AXI_05_RID;
    output AXI_05_RLAST;
    output [1:0] AXI_05_RRESP;
    output AXI_05_RVALID;
    output AXI_05_WREADY;
    output AXI_06_ARREADY;
    output AXI_06_AWREADY;
    output [5:0] AXI_06_BID;
    output [1:0] AXI_06_BRESP;
    output AXI_06_BVALID;
    output [1:0] AXI_06_DFI_AW_AERR_N;
    output AXI_06_DFI_CLK_BUF;
    output [7:0] AXI_06_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_06_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_06_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_06_DFI_DW_RDDATA_VALID;
    output AXI_06_DFI_INIT_COMPLETE;
    output AXI_06_DFI_PHYUPD_REQ;
    output AXI_06_DFI_PHY_LP_STATE;
    output AXI_06_DFI_RST_N_BUF;
    output [5:0] AXI_06_MC_STATUS;
    output [7:0] AXI_06_PHY_STATUS;
    output [255:0] AXI_06_RDATA;
    output [31:0] AXI_06_RDATA_PARITY;
    output [5:0] AXI_06_RID;
    output AXI_06_RLAST;
    output [1:0] AXI_06_RRESP;
    output AXI_06_RVALID;
    output AXI_06_WREADY;
    output AXI_07_ARREADY;
    output AXI_07_AWREADY;
    output [5:0] AXI_07_BID;
    output [1:0] AXI_07_BRESP;
    output AXI_07_BVALID;
    output [1:0] AXI_07_DFI_AW_AERR_N;
    output AXI_07_DFI_CLK_BUF;
    output [7:0] AXI_07_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_07_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_07_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_07_DFI_DW_RDDATA_VALID;
    output AXI_07_DFI_INIT_COMPLETE;
    output AXI_07_DFI_PHYUPD_REQ;
    output AXI_07_DFI_PHY_LP_STATE;
    output AXI_07_DFI_RST_N_BUF;
    output [255:0] AXI_07_RDATA;
    output [31:0] AXI_07_RDATA_PARITY;
    output [5:0] AXI_07_RID;
    output AXI_07_RLAST;
    output [1:0] AXI_07_RRESP;
    output AXI_07_RVALID;
    output AXI_07_WREADY;
    output AXI_08_ARREADY;
    output AXI_08_AWREADY;
    output [5:0] AXI_08_BID;
    output [1:0] AXI_08_BRESP;
    output AXI_08_BVALID;
    output [1:0] AXI_08_DFI_AW_AERR_N;
    output AXI_08_DFI_CLK_BUF;
    output [7:0] AXI_08_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_08_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_08_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_08_DFI_DW_RDDATA_VALID;
    output AXI_08_DFI_INIT_COMPLETE;
    output AXI_08_DFI_PHYUPD_REQ;
    output AXI_08_DFI_PHY_LP_STATE;
    output AXI_08_DFI_RST_N_BUF;
    output [5:0] AXI_08_MC_STATUS;
    output [7:0] AXI_08_PHY_STATUS;
    output [255:0] AXI_08_RDATA;
    output [31:0] AXI_08_RDATA_PARITY;
    output [5:0] AXI_08_RID;
    output AXI_08_RLAST;
    output [1:0] AXI_08_RRESP;
    output AXI_08_RVALID;
    output AXI_08_WREADY;
    output AXI_09_ARREADY;
    output AXI_09_AWREADY;
    output [5:0] AXI_09_BID;
    output [1:0] AXI_09_BRESP;
    output AXI_09_BVALID;
    output [1:0] AXI_09_DFI_AW_AERR_N;
    output AXI_09_DFI_CLK_BUF;
    output [7:0] AXI_09_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_09_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_09_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_09_DFI_DW_RDDATA_VALID;
    output AXI_09_DFI_INIT_COMPLETE;
    output AXI_09_DFI_PHYUPD_REQ;
    output AXI_09_DFI_PHY_LP_STATE;
    output AXI_09_DFI_RST_N_BUF;
    output [255:0] AXI_09_RDATA;
    output [31:0] AXI_09_RDATA_PARITY;
    output [5:0] AXI_09_RID;
    output AXI_09_RLAST;
    output [1:0] AXI_09_RRESP;
    output AXI_09_RVALID;
    output AXI_09_WREADY;
    output AXI_10_ARREADY;
    output AXI_10_AWREADY;
    output [5:0] AXI_10_BID;
    output [1:0] AXI_10_BRESP;
    output AXI_10_BVALID;
    output [1:0] AXI_10_DFI_AW_AERR_N;
    output AXI_10_DFI_CLK_BUF;
    output [7:0] AXI_10_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_10_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_10_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_10_DFI_DW_RDDATA_VALID;
    output AXI_10_DFI_INIT_COMPLETE;
    output AXI_10_DFI_PHYUPD_REQ;
    output AXI_10_DFI_PHY_LP_STATE;
    output AXI_10_DFI_RST_N_BUF;
    output [5:0] AXI_10_MC_STATUS;
    output [7:0] AXI_10_PHY_STATUS;
    output [255:0] AXI_10_RDATA;
    output [31:0] AXI_10_RDATA_PARITY;
    output [5:0] AXI_10_RID;
    output AXI_10_RLAST;
    output [1:0] AXI_10_RRESP;
    output AXI_10_RVALID;
    output AXI_10_WREADY;
    output AXI_11_ARREADY;
    output AXI_11_AWREADY;
    output [5:0] AXI_11_BID;
    output [1:0] AXI_11_BRESP;
    output AXI_11_BVALID;
    output [1:0] AXI_11_DFI_AW_AERR_N;
    output AXI_11_DFI_CLK_BUF;
    output [7:0] AXI_11_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_11_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_11_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_11_DFI_DW_RDDATA_VALID;
    output AXI_11_DFI_INIT_COMPLETE;
    output AXI_11_DFI_PHYUPD_REQ;
    output AXI_11_DFI_PHY_LP_STATE;
    output AXI_11_DFI_RST_N_BUF;
    output [255:0] AXI_11_RDATA;
    output [31:0] AXI_11_RDATA_PARITY;
    output [5:0] AXI_11_RID;
    output AXI_11_RLAST;
    output [1:0] AXI_11_RRESP;
    output AXI_11_RVALID;
    output AXI_11_WREADY;
    output AXI_12_ARREADY;
    output AXI_12_AWREADY;
    output [5:0] AXI_12_BID;
    output [1:0] AXI_12_BRESP;
    output AXI_12_BVALID;
    output [1:0] AXI_12_DFI_AW_AERR_N;
    output AXI_12_DFI_CLK_BUF;
    output [7:0] AXI_12_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_12_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_12_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_12_DFI_DW_RDDATA_VALID;
    output AXI_12_DFI_INIT_COMPLETE;
    output AXI_12_DFI_PHYUPD_REQ;
    output AXI_12_DFI_PHY_LP_STATE;
    output AXI_12_DFI_RST_N_BUF;
    output [5:0] AXI_12_MC_STATUS;
    output [7:0] AXI_12_PHY_STATUS;
    output [255:0] AXI_12_RDATA;
    output [31:0] AXI_12_RDATA_PARITY;
    output [5:0] AXI_12_RID;
    output AXI_12_RLAST;
    output [1:0] AXI_12_RRESP;
    output AXI_12_RVALID;
    output AXI_12_WREADY;
    output AXI_13_ARREADY;
    output AXI_13_AWREADY;
    output [5:0] AXI_13_BID;
    output [1:0] AXI_13_BRESP;
    output AXI_13_BVALID;
    output [1:0] AXI_13_DFI_AW_AERR_N;
    output AXI_13_DFI_CLK_BUF;
    output [7:0] AXI_13_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_13_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_13_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_13_DFI_DW_RDDATA_VALID;
    output AXI_13_DFI_INIT_COMPLETE;
    output AXI_13_DFI_PHYUPD_REQ;
    output AXI_13_DFI_PHY_LP_STATE;
    output AXI_13_DFI_RST_N_BUF;
    output [255:0] AXI_13_RDATA;
    output [31:0] AXI_13_RDATA_PARITY;
    output [5:0] AXI_13_RID;
    output AXI_13_RLAST;
    output [1:0] AXI_13_RRESP;
    output AXI_13_RVALID;
    output AXI_13_WREADY;
    output AXI_14_ARREADY;
    output AXI_14_AWREADY;
    output [5:0] AXI_14_BID;
    output [1:0] AXI_14_BRESP;
    output AXI_14_BVALID;
    output [1:0] AXI_14_DFI_AW_AERR_N;
    output AXI_14_DFI_CLK_BUF;
    output [7:0] AXI_14_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_14_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_14_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_14_DFI_DW_RDDATA_VALID;
    output AXI_14_DFI_INIT_COMPLETE;
    output AXI_14_DFI_PHYUPD_REQ;
    output AXI_14_DFI_PHY_LP_STATE;
    output AXI_14_DFI_RST_N_BUF;
    output [5:0] AXI_14_MC_STATUS;
    output [7:0] AXI_14_PHY_STATUS;
    output [255:0] AXI_14_RDATA;
    output [31:0] AXI_14_RDATA_PARITY;
    output [5:0] AXI_14_RID;
    output AXI_14_RLAST;
    output [1:0] AXI_14_RRESP;
    output AXI_14_RVALID;
    output AXI_14_WREADY;
    output AXI_15_ARREADY;
    output AXI_15_AWREADY;
    output [5:0] AXI_15_BID;
    output [1:0] AXI_15_BRESP;
    output AXI_15_BVALID;
    output [1:0] AXI_15_DFI_AW_AERR_N;
    output AXI_15_DFI_CLK_BUF;
    output [7:0] AXI_15_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_15_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_15_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_15_DFI_DW_RDDATA_VALID;
    output AXI_15_DFI_INIT_COMPLETE;
    output AXI_15_DFI_PHYUPD_REQ;
    output AXI_15_DFI_PHY_LP_STATE;
    output AXI_15_DFI_RST_N_BUF;
    output [255:0] AXI_15_RDATA;
    output [31:0] AXI_15_RDATA_PARITY;
    output [5:0] AXI_15_RID;
    output AXI_15_RLAST;
    output [1:0] AXI_15_RRESP;
    output AXI_15_RVALID;
    output AXI_15_WREADY;
    output DRAM_0_STAT_CATTRIP;
    output [2:0] DRAM_0_STAT_TEMP;
    input [21:0] APB_0_PADDR;
    (* invertible_pin = "IS_APB_0_PCLK_INVERTED" *)
    input APB_0_PCLK;
    input APB_0_PENABLE;
    (* invertible_pin = "IS_APB_0_PRESET_N_INVERTED" *)
    input APB_0_PRESET_N;
    input APB_0_PSEL;
    input [31:0] APB_0_PWDATA;
    input APB_0_PWRITE;
    (* invertible_pin = "IS_AXI_00_ACLK_INVERTED" *)
    input AXI_00_ACLK;
    input [36:0] AXI_00_ARADDR;
    input [1:0] AXI_00_ARBURST;
    (* invertible_pin = "IS_AXI_00_ARESET_N_INVERTED" *)
    input AXI_00_ARESET_N;
    input [5:0] AXI_00_ARID;
    input [3:0] AXI_00_ARLEN;
    input [2:0] AXI_00_ARSIZE;
    input AXI_00_ARVALID;
    input [36:0] AXI_00_AWADDR;
    input [1:0] AXI_00_AWBURST;
    input [5:0] AXI_00_AWID;
    input [3:0] AXI_00_AWLEN;
    input [2:0] AXI_00_AWSIZE;
    input AXI_00_AWVALID;
    input AXI_00_BREADY;
    input AXI_00_DFI_LP_PWR_X_REQ;
    input AXI_00_RREADY;
    input [255:0] AXI_00_WDATA;
    input [31:0] AXI_00_WDATA_PARITY;
    input AXI_00_WLAST;
    input [31:0] AXI_00_WSTRB;
    input AXI_00_WVALID;
    (* invertible_pin = "IS_AXI_01_ACLK_INVERTED" *)
    input AXI_01_ACLK;
    input [36:0] AXI_01_ARADDR;
    input [1:0] AXI_01_ARBURST;
    (* invertible_pin = "IS_AXI_01_ARESET_N_INVERTED" *)
    input AXI_01_ARESET_N;
    input [5:0] AXI_01_ARID;
    input [3:0] AXI_01_ARLEN;
    input [2:0] AXI_01_ARSIZE;
    input AXI_01_ARVALID;
    input [36:0] AXI_01_AWADDR;
    input [1:0] AXI_01_AWBURST;
    input [5:0] AXI_01_AWID;
    input [3:0] AXI_01_AWLEN;
    input [2:0] AXI_01_AWSIZE;
    input AXI_01_AWVALID;
    input AXI_01_BREADY;
    input AXI_01_DFI_LP_PWR_X_REQ;
    input AXI_01_RREADY;
    input [255:0] AXI_01_WDATA;
    input [31:0] AXI_01_WDATA_PARITY;
    input AXI_01_WLAST;
    input [31:0] AXI_01_WSTRB;
    input AXI_01_WVALID;
    (* invertible_pin = "IS_AXI_02_ACLK_INVERTED" *)
    input AXI_02_ACLK;
    input [36:0] AXI_02_ARADDR;
    input [1:0] AXI_02_ARBURST;
    (* invertible_pin = "IS_AXI_02_ARESET_N_INVERTED" *)
    input AXI_02_ARESET_N;
    input [5:0] AXI_02_ARID;
    input [3:0] AXI_02_ARLEN;
    input [2:0] AXI_02_ARSIZE;
    input AXI_02_ARVALID;
    input [36:0] AXI_02_AWADDR;
    input [1:0] AXI_02_AWBURST;
    input [5:0] AXI_02_AWID;
    input [3:0] AXI_02_AWLEN;
    input [2:0] AXI_02_AWSIZE;
    input AXI_02_AWVALID;
    input AXI_02_BREADY;
    input AXI_02_DFI_LP_PWR_X_REQ;
    input AXI_02_RREADY;
    input [255:0] AXI_02_WDATA;
    input [31:0] AXI_02_WDATA_PARITY;
    input AXI_02_WLAST;
    input [31:0] AXI_02_WSTRB;
    input AXI_02_WVALID;
    (* invertible_pin = "IS_AXI_03_ACLK_INVERTED" *)
    input AXI_03_ACLK;
    input [36:0] AXI_03_ARADDR;
    input [1:0] AXI_03_ARBURST;
    (* invertible_pin = "IS_AXI_03_ARESET_N_INVERTED" *)
    input AXI_03_ARESET_N;
    input [5:0] AXI_03_ARID;
    input [3:0] AXI_03_ARLEN;
    input [2:0] AXI_03_ARSIZE;
    input AXI_03_ARVALID;
    input [36:0] AXI_03_AWADDR;
    input [1:0] AXI_03_AWBURST;
    input [5:0] AXI_03_AWID;
    input [3:0] AXI_03_AWLEN;
    input [2:0] AXI_03_AWSIZE;
    input AXI_03_AWVALID;
    input AXI_03_BREADY;
    input AXI_03_DFI_LP_PWR_X_REQ;
    input AXI_03_RREADY;
    input [255:0] AXI_03_WDATA;
    input [31:0] AXI_03_WDATA_PARITY;
    input AXI_03_WLAST;
    input [31:0] AXI_03_WSTRB;
    input AXI_03_WVALID;
    (* invertible_pin = "IS_AXI_04_ACLK_INVERTED" *)
    input AXI_04_ACLK;
    input [36:0] AXI_04_ARADDR;
    input [1:0] AXI_04_ARBURST;
    (* invertible_pin = "IS_AXI_04_ARESET_N_INVERTED" *)
    input AXI_04_ARESET_N;
    input [5:0] AXI_04_ARID;
    input [3:0] AXI_04_ARLEN;
    input [2:0] AXI_04_ARSIZE;
    input AXI_04_ARVALID;
    input [36:0] AXI_04_AWADDR;
    input [1:0] AXI_04_AWBURST;
    input [5:0] AXI_04_AWID;
    input [3:0] AXI_04_AWLEN;
    input [2:0] AXI_04_AWSIZE;
    input AXI_04_AWVALID;
    input AXI_04_BREADY;
    input AXI_04_DFI_LP_PWR_X_REQ;
    input AXI_04_RREADY;
    input [255:0] AXI_04_WDATA;
    input [31:0] AXI_04_WDATA_PARITY;
    input AXI_04_WLAST;
    input [31:0] AXI_04_WSTRB;
    input AXI_04_WVALID;
    (* invertible_pin = "IS_AXI_05_ACLK_INVERTED" *)
    input AXI_05_ACLK;
    input [36:0] AXI_05_ARADDR;
    input [1:0] AXI_05_ARBURST;
    (* invertible_pin = "IS_AXI_05_ARESET_N_INVERTED" *)
    input AXI_05_ARESET_N;
    input [5:0] AXI_05_ARID;
    input [3:0] AXI_05_ARLEN;
    input [2:0] AXI_05_ARSIZE;
    input AXI_05_ARVALID;
    input [36:0] AXI_05_AWADDR;
    input [1:0] AXI_05_AWBURST;
    input [5:0] AXI_05_AWID;
    input [3:0] AXI_05_AWLEN;
    input [2:0] AXI_05_AWSIZE;
    input AXI_05_AWVALID;
    input AXI_05_BREADY;
    input AXI_05_DFI_LP_PWR_X_REQ;
    input AXI_05_RREADY;
    input [255:0] AXI_05_WDATA;
    input [31:0] AXI_05_WDATA_PARITY;
    input AXI_05_WLAST;
    input [31:0] AXI_05_WSTRB;
    input AXI_05_WVALID;
    (* invertible_pin = "IS_AXI_06_ACLK_INVERTED" *)
    input AXI_06_ACLK;
    input [36:0] AXI_06_ARADDR;
    input [1:0] AXI_06_ARBURST;
    (* invertible_pin = "IS_AXI_06_ARESET_N_INVERTED" *)
    input AXI_06_ARESET_N;
    input [5:0] AXI_06_ARID;
    input [3:0] AXI_06_ARLEN;
    input [2:0] AXI_06_ARSIZE;
    input AXI_06_ARVALID;
    input [36:0] AXI_06_AWADDR;
    input [1:0] AXI_06_AWBURST;
    input [5:0] AXI_06_AWID;
    input [3:0] AXI_06_AWLEN;
    input [2:0] AXI_06_AWSIZE;
    input AXI_06_AWVALID;
    input AXI_06_BREADY;
    input AXI_06_DFI_LP_PWR_X_REQ;
    input AXI_06_RREADY;
    input [255:0] AXI_06_WDATA;
    input [31:0] AXI_06_WDATA_PARITY;
    input AXI_06_WLAST;
    input [31:0] AXI_06_WSTRB;
    input AXI_06_WVALID;
    (* invertible_pin = "IS_AXI_07_ACLK_INVERTED" *)
    input AXI_07_ACLK;
    input [36:0] AXI_07_ARADDR;
    input [1:0] AXI_07_ARBURST;
    (* invertible_pin = "IS_AXI_07_ARESET_N_INVERTED" *)
    input AXI_07_ARESET_N;
    input [5:0] AXI_07_ARID;
    input [3:0] AXI_07_ARLEN;
    input [2:0] AXI_07_ARSIZE;
    input AXI_07_ARVALID;
    input [36:0] AXI_07_AWADDR;
    input [1:0] AXI_07_AWBURST;
    input [5:0] AXI_07_AWID;
    input [3:0] AXI_07_AWLEN;
    input [2:0] AXI_07_AWSIZE;
    input AXI_07_AWVALID;
    input AXI_07_BREADY;
    input AXI_07_DFI_LP_PWR_X_REQ;
    input AXI_07_RREADY;
    input [255:0] AXI_07_WDATA;
    input [31:0] AXI_07_WDATA_PARITY;
    input AXI_07_WLAST;
    input [31:0] AXI_07_WSTRB;
    input AXI_07_WVALID;
    (* invertible_pin = "IS_AXI_08_ACLK_INVERTED" *)
    input AXI_08_ACLK;
    input [36:0] AXI_08_ARADDR;
    input [1:0] AXI_08_ARBURST;
    (* invertible_pin = "IS_AXI_08_ARESET_N_INVERTED" *)
    input AXI_08_ARESET_N;
    input [5:0] AXI_08_ARID;
    input [3:0] AXI_08_ARLEN;
    input [2:0] AXI_08_ARSIZE;
    input AXI_08_ARVALID;
    input [36:0] AXI_08_AWADDR;
    input [1:0] AXI_08_AWBURST;
    input [5:0] AXI_08_AWID;
    input [3:0] AXI_08_AWLEN;
    input [2:0] AXI_08_AWSIZE;
    input AXI_08_AWVALID;
    input AXI_08_BREADY;
    input AXI_08_DFI_LP_PWR_X_REQ;
    input AXI_08_RREADY;
    input [255:0] AXI_08_WDATA;
    input [31:0] AXI_08_WDATA_PARITY;
    input AXI_08_WLAST;
    input [31:0] AXI_08_WSTRB;
    input AXI_08_WVALID;
    (* invertible_pin = "IS_AXI_09_ACLK_INVERTED" *)
    input AXI_09_ACLK;
    input [36:0] AXI_09_ARADDR;
    input [1:0] AXI_09_ARBURST;
    (* invertible_pin = "IS_AXI_09_ARESET_N_INVERTED" *)
    input AXI_09_ARESET_N;
    input [5:0] AXI_09_ARID;
    input [3:0] AXI_09_ARLEN;
    input [2:0] AXI_09_ARSIZE;
    input AXI_09_ARVALID;
    input [36:0] AXI_09_AWADDR;
    input [1:0] AXI_09_AWBURST;
    input [5:0] AXI_09_AWID;
    input [3:0] AXI_09_AWLEN;
    input [2:0] AXI_09_AWSIZE;
    input AXI_09_AWVALID;
    input AXI_09_BREADY;
    input AXI_09_DFI_LP_PWR_X_REQ;
    input AXI_09_RREADY;
    input [255:0] AXI_09_WDATA;
    input [31:0] AXI_09_WDATA_PARITY;
    input AXI_09_WLAST;
    input [31:0] AXI_09_WSTRB;
    input AXI_09_WVALID;
    (* invertible_pin = "IS_AXI_10_ACLK_INVERTED" *)
    input AXI_10_ACLK;
    input [36:0] AXI_10_ARADDR;
    input [1:0] AXI_10_ARBURST;
    (* invertible_pin = "IS_AXI_10_ARESET_N_INVERTED" *)
    input AXI_10_ARESET_N;
    input [5:0] AXI_10_ARID;
    input [3:0] AXI_10_ARLEN;
    input [2:0] AXI_10_ARSIZE;
    input AXI_10_ARVALID;
    input [36:0] AXI_10_AWADDR;
    input [1:0] AXI_10_AWBURST;
    input [5:0] AXI_10_AWID;
    input [3:0] AXI_10_AWLEN;
    input [2:0] AXI_10_AWSIZE;
    input AXI_10_AWVALID;
    input AXI_10_BREADY;
    input AXI_10_DFI_LP_PWR_X_REQ;
    input AXI_10_RREADY;
    input [255:0] AXI_10_WDATA;
    input [31:0] AXI_10_WDATA_PARITY;
    input AXI_10_WLAST;
    input [31:0] AXI_10_WSTRB;
    input AXI_10_WVALID;
    (* invertible_pin = "IS_AXI_11_ACLK_INVERTED" *)
    input AXI_11_ACLK;
    input [36:0] AXI_11_ARADDR;
    input [1:0] AXI_11_ARBURST;
    (* invertible_pin = "IS_AXI_11_ARESET_N_INVERTED" *)
    input AXI_11_ARESET_N;
    input [5:0] AXI_11_ARID;
    input [3:0] AXI_11_ARLEN;
    input [2:0] AXI_11_ARSIZE;
    input AXI_11_ARVALID;
    input [36:0] AXI_11_AWADDR;
    input [1:0] AXI_11_AWBURST;
    input [5:0] AXI_11_AWID;
    input [3:0] AXI_11_AWLEN;
    input [2:0] AXI_11_AWSIZE;
    input AXI_11_AWVALID;
    input AXI_11_BREADY;
    input AXI_11_DFI_LP_PWR_X_REQ;
    input AXI_11_RREADY;
    input [255:0] AXI_11_WDATA;
    input [31:0] AXI_11_WDATA_PARITY;
    input AXI_11_WLAST;
    input [31:0] AXI_11_WSTRB;
    input AXI_11_WVALID;
    (* invertible_pin = "IS_AXI_12_ACLK_INVERTED" *)
    input AXI_12_ACLK;
    input [36:0] AXI_12_ARADDR;
    input [1:0] AXI_12_ARBURST;
    (* invertible_pin = "IS_AXI_12_ARESET_N_INVERTED" *)
    input AXI_12_ARESET_N;
    input [5:0] AXI_12_ARID;
    input [3:0] AXI_12_ARLEN;
    input [2:0] AXI_12_ARSIZE;
    input AXI_12_ARVALID;
    input [36:0] AXI_12_AWADDR;
    input [1:0] AXI_12_AWBURST;
    input [5:0] AXI_12_AWID;
    input [3:0] AXI_12_AWLEN;
    input [2:0] AXI_12_AWSIZE;
    input AXI_12_AWVALID;
    input AXI_12_BREADY;
    input AXI_12_DFI_LP_PWR_X_REQ;
    input AXI_12_RREADY;
    input [255:0] AXI_12_WDATA;
    input [31:0] AXI_12_WDATA_PARITY;
    input AXI_12_WLAST;
    input [31:0] AXI_12_WSTRB;
    input AXI_12_WVALID;
    (* invertible_pin = "IS_AXI_13_ACLK_INVERTED" *)
    input AXI_13_ACLK;
    input [36:0] AXI_13_ARADDR;
    input [1:0] AXI_13_ARBURST;
    (* invertible_pin = "IS_AXI_13_ARESET_N_INVERTED" *)
    input AXI_13_ARESET_N;
    input [5:0] AXI_13_ARID;
    input [3:0] AXI_13_ARLEN;
    input [2:0] AXI_13_ARSIZE;
    input AXI_13_ARVALID;
    input [36:0] AXI_13_AWADDR;
    input [1:0] AXI_13_AWBURST;
    input [5:0] AXI_13_AWID;
    input [3:0] AXI_13_AWLEN;
    input [2:0] AXI_13_AWSIZE;
    input AXI_13_AWVALID;
    input AXI_13_BREADY;
    input AXI_13_DFI_LP_PWR_X_REQ;
    input AXI_13_RREADY;
    input [255:0] AXI_13_WDATA;
    input [31:0] AXI_13_WDATA_PARITY;
    input AXI_13_WLAST;
    input [31:0] AXI_13_WSTRB;
    input AXI_13_WVALID;
    (* invertible_pin = "IS_AXI_14_ACLK_INVERTED" *)
    input AXI_14_ACLK;
    input [36:0] AXI_14_ARADDR;
    input [1:0] AXI_14_ARBURST;
    (* invertible_pin = "IS_AXI_14_ARESET_N_INVERTED" *)
    input AXI_14_ARESET_N;
    input [5:0] AXI_14_ARID;
    input [3:0] AXI_14_ARLEN;
    input [2:0] AXI_14_ARSIZE;
    input AXI_14_ARVALID;
    input [36:0] AXI_14_AWADDR;
    input [1:0] AXI_14_AWBURST;
    input [5:0] AXI_14_AWID;
    input [3:0] AXI_14_AWLEN;
    input [2:0] AXI_14_AWSIZE;
    input AXI_14_AWVALID;
    input AXI_14_BREADY;
    input AXI_14_DFI_LP_PWR_X_REQ;
    input AXI_14_RREADY;
    input [255:0] AXI_14_WDATA;
    input [31:0] AXI_14_WDATA_PARITY;
    input AXI_14_WLAST;
    input [31:0] AXI_14_WSTRB;
    input AXI_14_WVALID;
    (* invertible_pin = "IS_AXI_15_ACLK_INVERTED" *)
    input AXI_15_ACLK;
    input [36:0] AXI_15_ARADDR;
    input [1:0] AXI_15_ARBURST;
    (* invertible_pin = "IS_AXI_15_ARESET_N_INVERTED" *)
    input AXI_15_ARESET_N;
    input [5:0] AXI_15_ARID;
    input [3:0] AXI_15_ARLEN;
    input [2:0] AXI_15_ARSIZE;
    input AXI_15_ARVALID;
    input [36:0] AXI_15_AWADDR;
    input [1:0] AXI_15_AWBURST;
    input [5:0] AXI_15_AWID;
    input [3:0] AXI_15_AWLEN;
    input [2:0] AXI_15_AWSIZE;
    input AXI_15_AWVALID;
    input AXI_15_BREADY;
    input AXI_15_DFI_LP_PWR_X_REQ;
    input AXI_15_RREADY;
    input [255:0] AXI_15_WDATA;
    input [31:0] AXI_15_WDATA_PARITY;
    input AXI_15_WLAST;
    input [31:0] AXI_15_WSTRB;
    input AXI_15_WVALID;
    input BSCAN_DRCK;
    input BSCAN_TCK;
    input HBM_REF_CLK;
    input MBIST_EN_00;
    input MBIST_EN_01;
    input MBIST_EN_02;
    input MBIST_EN_03;
    input MBIST_EN_04;
    input MBIST_EN_05;
    input MBIST_EN_06;
    input MBIST_EN_07;
endmodule

(* keep *)
module HBM_TWO_STACK_INTF (...);
    parameter CLK_SEL_00 = "FALSE";
    parameter CLK_SEL_01 = "FALSE";
    parameter CLK_SEL_02 = "FALSE";
    parameter CLK_SEL_03 = "FALSE";
    parameter CLK_SEL_04 = "FALSE";
    parameter CLK_SEL_05 = "FALSE";
    parameter CLK_SEL_06 = "FALSE";
    parameter CLK_SEL_07 = "FALSE";
    parameter CLK_SEL_08 = "FALSE";
    parameter CLK_SEL_09 = "FALSE";
    parameter CLK_SEL_10 = "FALSE";
    parameter CLK_SEL_11 = "FALSE";
    parameter CLK_SEL_12 = "FALSE";
    parameter CLK_SEL_13 = "FALSE";
    parameter CLK_SEL_14 = "FALSE";
    parameter CLK_SEL_15 = "FALSE";
    parameter CLK_SEL_16 = "FALSE";
    parameter CLK_SEL_17 = "FALSE";
    parameter CLK_SEL_18 = "FALSE";
    parameter CLK_SEL_19 = "FALSE";
    parameter CLK_SEL_20 = "FALSE";
    parameter CLK_SEL_21 = "FALSE";
    parameter CLK_SEL_22 = "FALSE";
    parameter CLK_SEL_23 = "FALSE";
    parameter CLK_SEL_24 = "FALSE";
    parameter CLK_SEL_25 = "FALSE";
    parameter CLK_SEL_26 = "FALSE";
    parameter CLK_SEL_27 = "FALSE";
    parameter CLK_SEL_28 = "FALSE";
    parameter CLK_SEL_29 = "FALSE";
    parameter CLK_SEL_30 = "FALSE";
    parameter CLK_SEL_31 = "FALSE";
    parameter integer DATARATE_00 = 1800;
    parameter integer DATARATE_01 = 1800;
    parameter integer DATARATE_02 = 1800;
    parameter integer DATARATE_03 = 1800;
    parameter integer DATARATE_04 = 1800;
    parameter integer DATARATE_05 = 1800;
    parameter integer DATARATE_06 = 1800;
    parameter integer DATARATE_07 = 1800;
    parameter integer DATARATE_08 = 1800;
    parameter integer DATARATE_09 = 1800;
    parameter integer DATARATE_10 = 1800;
    parameter integer DATARATE_11 = 1800;
    parameter integer DATARATE_12 = 1800;
    parameter integer DATARATE_13 = 1800;
    parameter integer DATARATE_14 = 1800;
    parameter integer DATARATE_15 = 1800;
    parameter DA_LOCKOUT_0 = "FALSE";
    parameter DA_LOCKOUT_1 = "FALSE";
    parameter [0:0] IS_APB_0_PCLK_INVERTED = 1'b0;
    parameter [0:0] IS_APB_0_PRESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_APB_1_PCLK_INVERTED = 1'b0;
    parameter [0:0] IS_APB_1_PRESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_00_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_00_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_01_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_01_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_02_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_02_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_03_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_03_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_04_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_04_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_05_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_05_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_06_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_06_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_07_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_07_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_08_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_08_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_09_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_09_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_10_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_10_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_11_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_11_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_12_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_12_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_13_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_13_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_14_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_14_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_15_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_15_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_16_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_16_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_17_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_17_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_18_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_18_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_19_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_19_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_20_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_20_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_21_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_21_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_22_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_22_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_23_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_23_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_24_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_24_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_25_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_25_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_26_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_26_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_27_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_27_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_28_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_28_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_29_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_29_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_30_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_30_ARESET_N_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_31_ACLK_INVERTED = 1'b0;
    parameter [0:0] IS_AXI_31_ARESET_N_INVERTED = 1'b0;
    parameter MC_ENABLE_00 = "FALSE";
    parameter MC_ENABLE_01 = "FALSE";
    parameter MC_ENABLE_02 = "FALSE";
    parameter MC_ENABLE_03 = "FALSE";
    parameter MC_ENABLE_04 = "FALSE";
    parameter MC_ENABLE_05 = "FALSE";
    parameter MC_ENABLE_06 = "FALSE";
    parameter MC_ENABLE_07 = "FALSE";
    parameter MC_ENABLE_08 = "FALSE";
    parameter MC_ENABLE_09 = "FALSE";
    parameter MC_ENABLE_10 = "FALSE";
    parameter MC_ENABLE_11 = "FALSE";
    parameter MC_ENABLE_12 = "FALSE";
    parameter MC_ENABLE_13 = "FALSE";
    parameter MC_ENABLE_14 = "FALSE";
    parameter MC_ENABLE_15 = "FALSE";
    parameter MC_ENABLE_APB_00 = "FALSE";
    parameter MC_ENABLE_APB_01 = "FALSE";
    parameter integer PAGEHIT_PERCENT_00 = 75;
    parameter integer PAGEHIT_PERCENT_01 = 75;
    parameter PHY_ENABLE_00 = "FALSE";
    parameter PHY_ENABLE_01 = "FALSE";
    parameter PHY_ENABLE_02 = "FALSE";
    parameter PHY_ENABLE_03 = "FALSE";
    parameter PHY_ENABLE_04 = "FALSE";
    parameter PHY_ENABLE_05 = "FALSE";
    parameter PHY_ENABLE_06 = "FALSE";
    parameter PHY_ENABLE_07 = "FALSE";
    parameter PHY_ENABLE_08 = "FALSE";
    parameter PHY_ENABLE_09 = "FALSE";
    parameter PHY_ENABLE_10 = "FALSE";
    parameter PHY_ENABLE_11 = "FALSE";
    parameter PHY_ENABLE_12 = "FALSE";
    parameter PHY_ENABLE_13 = "FALSE";
    parameter PHY_ENABLE_14 = "FALSE";
    parameter PHY_ENABLE_15 = "FALSE";
    parameter PHY_ENABLE_16 = "FALSE";
    parameter PHY_ENABLE_17 = "FALSE";
    parameter PHY_ENABLE_18 = "FALSE";
    parameter PHY_ENABLE_19 = "FALSE";
    parameter PHY_ENABLE_20 = "FALSE";
    parameter PHY_ENABLE_21 = "FALSE";
    parameter PHY_ENABLE_22 = "FALSE";
    parameter PHY_ENABLE_23 = "FALSE";
    parameter PHY_ENABLE_24 = "FALSE";
    parameter PHY_ENABLE_25 = "FALSE";
    parameter PHY_ENABLE_26 = "FALSE";
    parameter PHY_ENABLE_27 = "FALSE";
    parameter PHY_ENABLE_28 = "FALSE";
    parameter PHY_ENABLE_29 = "FALSE";
    parameter PHY_ENABLE_30 = "FALSE";
    parameter PHY_ENABLE_31 = "FALSE";
    parameter PHY_ENABLE_APB_00 = "FALSE";
    parameter PHY_ENABLE_APB_01 = "FALSE";
    parameter PHY_PCLK_INVERT_01 = "FALSE";
    parameter PHY_PCLK_INVERT_02 = "FALSE";
    parameter integer READ_PERCENT_00 = 50;
    parameter integer READ_PERCENT_01 = 50;
    parameter integer READ_PERCENT_02 = 50;
    parameter integer READ_PERCENT_03 = 50;
    parameter integer READ_PERCENT_04 = 50;
    parameter integer READ_PERCENT_05 = 50;
    parameter integer READ_PERCENT_06 = 50;
    parameter integer READ_PERCENT_07 = 50;
    parameter integer READ_PERCENT_08 = 50;
    parameter integer READ_PERCENT_09 = 50;
    parameter integer READ_PERCENT_10 = 50;
    parameter integer READ_PERCENT_11 = 50;
    parameter integer READ_PERCENT_12 = 50;
    parameter integer READ_PERCENT_13 = 50;
    parameter integer READ_PERCENT_14 = 50;
    parameter integer READ_PERCENT_15 = 50;
    parameter integer READ_PERCENT_16 = 50;
    parameter integer READ_PERCENT_17 = 50;
    parameter integer READ_PERCENT_18 = 50;
    parameter integer READ_PERCENT_19 = 50;
    parameter integer READ_PERCENT_20 = 50;
    parameter integer READ_PERCENT_21 = 50;
    parameter integer READ_PERCENT_22 = 50;
    parameter integer READ_PERCENT_23 = 50;
    parameter integer READ_PERCENT_24 = 50;
    parameter integer READ_PERCENT_25 = 50;
    parameter integer READ_PERCENT_26 = 50;
    parameter integer READ_PERCENT_27 = 50;
    parameter integer READ_PERCENT_28 = 50;
    parameter integer READ_PERCENT_29 = 50;
    parameter integer READ_PERCENT_30 = 50;
    parameter integer READ_PERCENT_31 = 50;
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter SWITCH_ENABLE_00 = "FALSE";
    parameter SWITCH_ENABLE_01 = "FALSE";
    parameter integer WRITE_PERCENT_00 = 50;
    parameter integer WRITE_PERCENT_01 = 50;
    parameter integer WRITE_PERCENT_02 = 50;
    parameter integer WRITE_PERCENT_03 = 50;
    parameter integer WRITE_PERCENT_04 = 50;
    parameter integer WRITE_PERCENT_05 = 50;
    parameter integer WRITE_PERCENT_06 = 50;
    parameter integer WRITE_PERCENT_07 = 50;
    parameter integer WRITE_PERCENT_08 = 50;
    parameter integer WRITE_PERCENT_09 = 50;
    parameter integer WRITE_PERCENT_10 = 50;
    parameter integer WRITE_PERCENT_11 = 50;
    parameter integer WRITE_PERCENT_12 = 50;
    parameter integer WRITE_PERCENT_13 = 50;
    parameter integer WRITE_PERCENT_14 = 50;
    parameter integer WRITE_PERCENT_15 = 50;
    parameter integer WRITE_PERCENT_16 = 50;
    parameter integer WRITE_PERCENT_17 = 50;
    parameter integer WRITE_PERCENT_18 = 50;
    parameter integer WRITE_PERCENT_19 = 50;
    parameter integer WRITE_PERCENT_20 = 50;
    parameter integer WRITE_PERCENT_21 = 50;
    parameter integer WRITE_PERCENT_22 = 50;
    parameter integer WRITE_PERCENT_23 = 50;
    parameter integer WRITE_PERCENT_24 = 50;
    parameter integer WRITE_PERCENT_25 = 50;
    parameter integer WRITE_PERCENT_26 = 50;
    parameter integer WRITE_PERCENT_27 = 50;
    parameter integer WRITE_PERCENT_28 = 50;
    parameter integer WRITE_PERCENT_29 = 50;
    parameter integer WRITE_PERCENT_30 = 50;
    parameter integer WRITE_PERCENT_31 = 50;
    output [31:0] APB_0_PRDATA;
    output APB_0_PREADY;
    output APB_0_PSLVERR;
    output [31:0] APB_1_PRDATA;
    output APB_1_PREADY;
    output APB_1_PSLVERR;
    output AXI_00_ARREADY;
    output AXI_00_AWREADY;
    output [5:0] AXI_00_BID;
    output [1:0] AXI_00_BRESP;
    output AXI_00_BVALID;
    output [1:0] AXI_00_DFI_AW_AERR_N;
    output AXI_00_DFI_CLK_BUF;
    output [7:0] AXI_00_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_00_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_00_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_00_DFI_DW_RDDATA_VALID;
    output AXI_00_DFI_INIT_COMPLETE;
    output AXI_00_DFI_PHYUPD_REQ;
    output AXI_00_DFI_PHY_LP_STATE;
    output AXI_00_DFI_RST_N_BUF;
    output [5:0] AXI_00_MC_STATUS;
    output [7:0] AXI_00_PHY_STATUS;
    output [255:0] AXI_00_RDATA;
    output [31:0] AXI_00_RDATA_PARITY;
    output [5:0] AXI_00_RID;
    output AXI_00_RLAST;
    output [1:0] AXI_00_RRESP;
    output AXI_00_RVALID;
    output AXI_00_WREADY;
    output AXI_01_ARREADY;
    output AXI_01_AWREADY;
    output [5:0] AXI_01_BID;
    output [1:0] AXI_01_BRESP;
    output AXI_01_BVALID;
    output [1:0] AXI_01_DFI_AW_AERR_N;
    output AXI_01_DFI_CLK_BUF;
    output [7:0] AXI_01_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_01_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_01_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_01_DFI_DW_RDDATA_VALID;
    output AXI_01_DFI_INIT_COMPLETE;
    output AXI_01_DFI_PHYUPD_REQ;
    output AXI_01_DFI_PHY_LP_STATE;
    output AXI_01_DFI_RST_N_BUF;
    output [255:0] AXI_01_RDATA;
    output [31:0] AXI_01_RDATA_PARITY;
    output [5:0] AXI_01_RID;
    output AXI_01_RLAST;
    output [1:0] AXI_01_RRESP;
    output AXI_01_RVALID;
    output AXI_01_WREADY;
    output AXI_02_ARREADY;
    output AXI_02_AWREADY;
    output [5:0] AXI_02_BID;
    output [1:0] AXI_02_BRESP;
    output AXI_02_BVALID;
    output [1:0] AXI_02_DFI_AW_AERR_N;
    output AXI_02_DFI_CLK_BUF;
    output [7:0] AXI_02_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_02_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_02_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_02_DFI_DW_RDDATA_VALID;
    output AXI_02_DFI_INIT_COMPLETE;
    output AXI_02_DFI_PHYUPD_REQ;
    output AXI_02_DFI_PHY_LP_STATE;
    output AXI_02_DFI_RST_N_BUF;
    output [5:0] AXI_02_MC_STATUS;
    output [7:0] AXI_02_PHY_STATUS;
    output [255:0] AXI_02_RDATA;
    output [31:0] AXI_02_RDATA_PARITY;
    output [5:0] AXI_02_RID;
    output AXI_02_RLAST;
    output [1:0] AXI_02_RRESP;
    output AXI_02_RVALID;
    output AXI_02_WREADY;
    output AXI_03_ARREADY;
    output AXI_03_AWREADY;
    output [5:0] AXI_03_BID;
    output [1:0] AXI_03_BRESP;
    output AXI_03_BVALID;
    output [1:0] AXI_03_DFI_AW_AERR_N;
    output AXI_03_DFI_CLK_BUF;
    output [7:0] AXI_03_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_03_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_03_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_03_DFI_DW_RDDATA_VALID;
    output AXI_03_DFI_INIT_COMPLETE;
    output AXI_03_DFI_PHYUPD_REQ;
    output AXI_03_DFI_PHY_LP_STATE;
    output AXI_03_DFI_RST_N_BUF;
    output [255:0] AXI_03_RDATA;
    output [31:0] AXI_03_RDATA_PARITY;
    output [5:0] AXI_03_RID;
    output AXI_03_RLAST;
    output [1:0] AXI_03_RRESP;
    output AXI_03_RVALID;
    output AXI_03_WREADY;
    output AXI_04_ARREADY;
    output AXI_04_AWREADY;
    output [5:0] AXI_04_BID;
    output [1:0] AXI_04_BRESP;
    output AXI_04_BVALID;
    output [1:0] AXI_04_DFI_AW_AERR_N;
    output AXI_04_DFI_CLK_BUF;
    output [7:0] AXI_04_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_04_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_04_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_04_DFI_DW_RDDATA_VALID;
    output AXI_04_DFI_INIT_COMPLETE;
    output AXI_04_DFI_PHYUPD_REQ;
    output AXI_04_DFI_PHY_LP_STATE;
    output AXI_04_DFI_RST_N_BUF;
    output [5:0] AXI_04_MC_STATUS;
    output [7:0] AXI_04_PHY_STATUS;
    output [255:0] AXI_04_RDATA;
    output [31:0] AXI_04_RDATA_PARITY;
    output [5:0] AXI_04_RID;
    output AXI_04_RLAST;
    output [1:0] AXI_04_RRESP;
    output AXI_04_RVALID;
    output AXI_04_WREADY;
    output AXI_05_ARREADY;
    output AXI_05_AWREADY;
    output [5:0] AXI_05_BID;
    output [1:0] AXI_05_BRESP;
    output AXI_05_BVALID;
    output [1:0] AXI_05_DFI_AW_AERR_N;
    output AXI_05_DFI_CLK_BUF;
    output [7:0] AXI_05_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_05_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_05_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_05_DFI_DW_RDDATA_VALID;
    output AXI_05_DFI_INIT_COMPLETE;
    output AXI_05_DFI_PHYUPD_REQ;
    output AXI_05_DFI_PHY_LP_STATE;
    output AXI_05_DFI_RST_N_BUF;
    output [255:0] AXI_05_RDATA;
    output [31:0] AXI_05_RDATA_PARITY;
    output [5:0] AXI_05_RID;
    output AXI_05_RLAST;
    output [1:0] AXI_05_RRESP;
    output AXI_05_RVALID;
    output AXI_05_WREADY;
    output AXI_06_ARREADY;
    output AXI_06_AWREADY;
    output [5:0] AXI_06_BID;
    output [1:0] AXI_06_BRESP;
    output AXI_06_BVALID;
    output [1:0] AXI_06_DFI_AW_AERR_N;
    output AXI_06_DFI_CLK_BUF;
    output [7:0] AXI_06_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_06_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_06_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_06_DFI_DW_RDDATA_VALID;
    output AXI_06_DFI_INIT_COMPLETE;
    output AXI_06_DFI_PHYUPD_REQ;
    output AXI_06_DFI_PHY_LP_STATE;
    output AXI_06_DFI_RST_N_BUF;
    output [5:0] AXI_06_MC_STATUS;
    output [7:0] AXI_06_PHY_STATUS;
    output [255:0] AXI_06_RDATA;
    output [31:0] AXI_06_RDATA_PARITY;
    output [5:0] AXI_06_RID;
    output AXI_06_RLAST;
    output [1:0] AXI_06_RRESP;
    output AXI_06_RVALID;
    output AXI_06_WREADY;
    output AXI_07_ARREADY;
    output AXI_07_AWREADY;
    output [5:0] AXI_07_BID;
    output [1:0] AXI_07_BRESP;
    output AXI_07_BVALID;
    output [1:0] AXI_07_DFI_AW_AERR_N;
    output AXI_07_DFI_CLK_BUF;
    output [7:0] AXI_07_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_07_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_07_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_07_DFI_DW_RDDATA_VALID;
    output AXI_07_DFI_INIT_COMPLETE;
    output AXI_07_DFI_PHYUPD_REQ;
    output AXI_07_DFI_PHY_LP_STATE;
    output AXI_07_DFI_RST_N_BUF;
    output [255:0] AXI_07_RDATA;
    output [31:0] AXI_07_RDATA_PARITY;
    output [5:0] AXI_07_RID;
    output AXI_07_RLAST;
    output [1:0] AXI_07_RRESP;
    output AXI_07_RVALID;
    output AXI_07_WREADY;
    output AXI_08_ARREADY;
    output AXI_08_AWREADY;
    output [5:0] AXI_08_BID;
    output [1:0] AXI_08_BRESP;
    output AXI_08_BVALID;
    output [1:0] AXI_08_DFI_AW_AERR_N;
    output AXI_08_DFI_CLK_BUF;
    output [7:0] AXI_08_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_08_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_08_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_08_DFI_DW_RDDATA_VALID;
    output AXI_08_DFI_INIT_COMPLETE;
    output AXI_08_DFI_PHYUPD_REQ;
    output AXI_08_DFI_PHY_LP_STATE;
    output AXI_08_DFI_RST_N_BUF;
    output [5:0] AXI_08_MC_STATUS;
    output [7:0] AXI_08_PHY_STATUS;
    output [255:0] AXI_08_RDATA;
    output [31:0] AXI_08_RDATA_PARITY;
    output [5:0] AXI_08_RID;
    output AXI_08_RLAST;
    output [1:0] AXI_08_RRESP;
    output AXI_08_RVALID;
    output AXI_08_WREADY;
    output AXI_09_ARREADY;
    output AXI_09_AWREADY;
    output [5:0] AXI_09_BID;
    output [1:0] AXI_09_BRESP;
    output AXI_09_BVALID;
    output [1:0] AXI_09_DFI_AW_AERR_N;
    output AXI_09_DFI_CLK_BUF;
    output [7:0] AXI_09_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_09_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_09_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_09_DFI_DW_RDDATA_VALID;
    output AXI_09_DFI_INIT_COMPLETE;
    output AXI_09_DFI_PHYUPD_REQ;
    output AXI_09_DFI_PHY_LP_STATE;
    output AXI_09_DFI_RST_N_BUF;
    output [255:0] AXI_09_RDATA;
    output [31:0] AXI_09_RDATA_PARITY;
    output [5:0] AXI_09_RID;
    output AXI_09_RLAST;
    output [1:0] AXI_09_RRESP;
    output AXI_09_RVALID;
    output AXI_09_WREADY;
    output AXI_10_ARREADY;
    output AXI_10_AWREADY;
    output [5:0] AXI_10_BID;
    output [1:0] AXI_10_BRESP;
    output AXI_10_BVALID;
    output [1:0] AXI_10_DFI_AW_AERR_N;
    output AXI_10_DFI_CLK_BUF;
    output [7:0] AXI_10_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_10_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_10_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_10_DFI_DW_RDDATA_VALID;
    output AXI_10_DFI_INIT_COMPLETE;
    output AXI_10_DFI_PHYUPD_REQ;
    output AXI_10_DFI_PHY_LP_STATE;
    output AXI_10_DFI_RST_N_BUF;
    output [5:0] AXI_10_MC_STATUS;
    output [7:0] AXI_10_PHY_STATUS;
    output [255:0] AXI_10_RDATA;
    output [31:0] AXI_10_RDATA_PARITY;
    output [5:0] AXI_10_RID;
    output AXI_10_RLAST;
    output [1:0] AXI_10_RRESP;
    output AXI_10_RVALID;
    output AXI_10_WREADY;
    output AXI_11_ARREADY;
    output AXI_11_AWREADY;
    output [5:0] AXI_11_BID;
    output [1:0] AXI_11_BRESP;
    output AXI_11_BVALID;
    output [1:0] AXI_11_DFI_AW_AERR_N;
    output AXI_11_DFI_CLK_BUF;
    output [7:0] AXI_11_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_11_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_11_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_11_DFI_DW_RDDATA_VALID;
    output AXI_11_DFI_INIT_COMPLETE;
    output AXI_11_DFI_PHYUPD_REQ;
    output AXI_11_DFI_PHY_LP_STATE;
    output AXI_11_DFI_RST_N_BUF;
    output [255:0] AXI_11_RDATA;
    output [31:0] AXI_11_RDATA_PARITY;
    output [5:0] AXI_11_RID;
    output AXI_11_RLAST;
    output [1:0] AXI_11_RRESP;
    output AXI_11_RVALID;
    output AXI_11_WREADY;
    output AXI_12_ARREADY;
    output AXI_12_AWREADY;
    output [5:0] AXI_12_BID;
    output [1:0] AXI_12_BRESP;
    output AXI_12_BVALID;
    output [1:0] AXI_12_DFI_AW_AERR_N;
    output AXI_12_DFI_CLK_BUF;
    output [7:0] AXI_12_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_12_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_12_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_12_DFI_DW_RDDATA_VALID;
    output AXI_12_DFI_INIT_COMPLETE;
    output AXI_12_DFI_PHYUPD_REQ;
    output AXI_12_DFI_PHY_LP_STATE;
    output AXI_12_DFI_RST_N_BUF;
    output [5:0] AXI_12_MC_STATUS;
    output [7:0] AXI_12_PHY_STATUS;
    output [255:0] AXI_12_RDATA;
    output [31:0] AXI_12_RDATA_PARITY;
    output [5:0] AXI_12_RID;
    output AXI_12_RLAST;
    output [1:0] AXI_12_RRESP;
    output AXI_12_RVALID;
    output AXI_12_WREADY;
    output AXI_13_ARREADY;
    output AXI_13_AWREADY;
    output [5:0] AXI_13_BID;
    output [1:0] AXI_13_BRESP;
    output AXI_13_BVALID;
    output [1:0] AXI_13_DFI_AW_AERR_N;
    output AXI_13_DFI_CLK_BUF;
    output [7:0] AXI_13_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_13_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_13_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_13_DFI_DW_RDDATA_VALID;
    output AXI_13_DFI_INIT_COMPLETE;
    output AXI_13_DFI_PHYUPD_REQ;
    output AXI_13_DFI_PHY_LP_STATE;
    output AXI_13_DFI_RST_N_BUF;
    output [255:0] AXI_13_RDATA;
    output [31:0] AXI_13_RDATA_PARITY;
    output [5:0] AXI_13_RID;
    output AXI_13_RLAST;
    output [1:0] AXI_13_RRESP;
    output AXI_13_RVALID;
    output AXI_13_WREADY;
    output AXI_14_ARREADY;
    output AXI_14_AWREADY;
    output [5:0] AXI_14_BID;
    output [1:0] AXI_14_BRESP;
    output AXI_14_BVALID;
    output [1:0] AXI_14_DFI_AW_AERR_N;
    output AXI_14_DFI_CLK_BUF;
    output [7:0] AXI_14_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_14_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_14_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_14_DFI_DW_RDDATA_VALID;
    output AXI_14_DFI_INIT_COMPLETE;
    output AXI_14_DFI_PHYUPD_REQ;
    output AXI_14_DFI_PHY_LP_STATE;
    output AXI_14_DFI_RST_N_BUF;
    output [5:0] AXI_14_MC_STATUS;
    output [7:0] AXI_14_PHY_STATUS;
    output [255:0] AXI_14_RDATA;
    output [31:0] AXI_14_RDATA_PARITY;
    output [5:0] AXI_14_RID;
    output AXI_14_RLAST;
    output [1:0] AXI_14_RRESP;
    output AXI_14_RVALID;
    output AXI_14_WREADY;
    output AXI_15_ARREADY;
    output AXI_15_AWREADY;
    output [5:0] AXI_15_BID;
    output [1:0] AXI_15_BRESP;
    output AXI_15_BVALID;
    output [1:0] AXI_15_DFI_AW_AERR_N;
    output AXI_15_DFI_CLK_BUF;
    output [7:0] AXI_15_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_15_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_15_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_15_DFI_DW_RDDATA_VALID;
    output AXI_15_DFI_INIT_COMPLETE;
    output AXI_15_DFI_PHYUPD_REQ;
    output AXI_15_DFI_PHY_LP_STATE;
    output AXI_15_DFI_RST_N_BUF;
    output [255:0] AXI_15_RDATA;
    output [31:0] AXI_15_RDATA_PARITY;
    output [5:0] AXI_15_RID;
    output AXI_15_RLAST;
    output [1:0] AXI_15_RRESP;
    output AXI_15_RVALID;
    output AXI_15_WREADY;
    output AXI_16_ARREADY;
    output AXI_16_AWREADY;
    output [5:0] AXI_16_BID;
    output [1:0] AXI_16_BRESP;
    output AXI_16_BVALID;
    output [1:0] AXI_16_DFI_AW_AERR_N;
    output AXI_16_DFI_CLK_BUF;
    output [7:0] AXI_16_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_16_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_16_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_16_DFI_DW_RDDATA_VALID;
    output AXI_16_DFI_INIT_COMPLETE;
    output AXI_16_DFI_PHYUPD_REQ;
    output AXI_16_DFI_PHY_LP_STATE;
    output AXI_16_DFI_RST_N_BUF;
    output [5:0] AXI_16_MC_STATUS;
    output [7:0] AXI_16_PHY_STATUS;
    output [255:0] AXI_16_RDATA;
    output [31:0] AXI_16_RDATA_PARITY;
    output [5:0] AXI_16_RID;
    output AXI_16_RLAST;
    output [1:0] AXI_16_RRESP;
    output AXI_16_RVALID;
    output AXI_16_WREADY;
    output AXI_17_ARREADY;
    output AXI_17_AWREADY;
    output [5:0] AXI_17_BID;
    output [1:0] AXI_17_BRESP;
    output AXI_17_BVALID;
    output [1:0] AXI_17_DFI_AW_AERR_N;
    output AXI_17_DFI_CLK_BUF;
    output [7:0] AXI_17_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_17_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_17_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_17_DFI_DW_RDDATA_VALID;
    output AXI_17_DFI_INIT_COMPLETE;
    output AXI_17_DFI_PHYUPD_REQ;
    output AXI_17_DFI_PHY_LP_STATE;
    output AXI_17_DFI_RST_N_BUF;
    output [255:0] AXI_17_RDATA;
    output [31:0] AXI_17_RDATA_PARITY;
    output [5:0] AXI_17_RID;
    output AXI_17_RLAST;
    output [1:0] AXI_17_RRESP;
    output AXI_17_RVALID;
    output AXI_17_WREADY;
    output AXI_18_ARREADY;
    output AXI_18_AWREADY;
    output [5:0] AXI_18_BID;
    output [1:0] AXI_18_BRESP;
    output AXI_18_BVALID;
    output [1:0] AXI_18_DFI_AW_AERR_N;
    output AXI_18_DFI_CLK_BUF;
    output [7:0] AXI_18_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_18_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_18_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_18_DFI_DW_RDDATA_VALID;
    output AXI_18_DFI_INIT_COMPLETE;
    output AXI_18_DFI_PHYUPD_REQ;
    output AXI_18_DFI_PHY_LP_STATE;
    output AXI_18_DFI_RST_N_BUF;
    output [5:0] AXI_18_MC_STATUS;
    output [7:0] AXI_18_PHY_STATUS;
    output [255:0] AXI_18_RDATA;
    output [31:0] AXI_18_RDATA_PARITY;
    output [5:0] AXI_18_RID;
    output AXI_18_RLAST;
    output [1:0] AXI_18_RRESP;
    output AXI_18_RVALID;
    output AXI_18_WREADY;
    output AXI_19_ARREADY;
    output AXI_19_AWREADY;
    output [5:0] AXI_19_BID;
    output [1:0] AXI_19_BRESP;
    output AXI_19_BVALID;
    output [1:0] AXI_19_DFI_AW_AERR_N;
    output AXI_19_DFI_CLK_BUF;
    output [7:0] AXI_19_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_19_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_19_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_19_DFI_DW_RDDATA_VALID;
    output AXI_19_DFI_INIT_COMPLETE;
    output AXI_19_DFI_PHYUPD_REQ;
    output AXI_19_DFI_PHY_LP_STATE;
    output AXI_19_DFI_RST_N_BUF;
    output [255:0] AXI_19_RDATA;
    output [31:0] AXI_19_RDATA_PARITY;
    output [5:0] AXI_19_RID;
    output AXI_19_RLAST;
    output [1:0] AXI_19_RRESP;
    output AXI_19_RVALID;
    output AXI_19_WREADY;
    output AXI_20_ARREADY;
    output AXI_20_AWREADY;
    output [5:0] AXI_20_BID;
    output [1:0] AXI_20_BRESP;
    output AXI_20_BVALID;
    output [1:0] AXI_20_DFI_AW_AERR_N;
    output AXI_20_DFI_CLK_BUF;
    output [7:0] AXI_20_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_20_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_20_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_20_DFI_DW_RDDATA_VALID;
    output AXI_20_DFI_INIT_COMPLETE;
    output AXI_20_DFI_PHYUPD_REQ;
    output AXI_20_DFI_PHY_LP_STATE;
    output AXI_20_DFI_RST_N_BUF;
    output [5:0] AXI_20_MC_STATUS;
    output [7:0] AXI_20_PHY_STATUS;
    output [255:0] AXI_20_RDATA;
    output [31:0] AXI_20_RDATA_PARITY;
    output [5:0] AXI_20_RID;
    output AXI_20_RLAST;
    output [1:0] AXI_20_RRESP;
    output AXI_20_RVALID;
    output AXI_20_WREADY;
    output AXI_21_ARREADY;
    output AXI_21_AWREADY;
    output [5:0] AXI_21_BID;
    output [1:0] AXI_21_BRESP;
    output AXI_21_BVALID;
    output [1:0] AXI_21_DFI_AW_AERR_N;
    output AXI_21_DFI_CLK_BUF;
    output [7:0] AXI_21_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_21_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_21_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_21_DFI_DW_RDDATA_VALID;
    output AXI_21_DFI_INIT_COMPLETE;
    output AXI_21_DFI_PHYUPD_REQ;
    output AXI_21_DFI_PHY_LP_STATE;
    output AXI_21_DFI_RST_N_BUF;
    output [255:0] AXI_21_RDATA;
    output [31:0] AXI_21_RDATA_PARITY;
    output [5:0] AXI_21_RID;
    output AXI_21_RLAST;
    output [1:0] AXI_21_RRESP;
    output AXI_21_RVALID;
    output AXI_21_WREADY;
    output AXI_22_ARREADY;
    output AXI_22_AWREADY;
    output [5:0] AXI_22_BID;
    output [1:0] AXI_22_BRESP;
    output AXI_22_BVALID;
    output [1:0] AXI_22_DFI_AW_AERR_N;
    output AXI_22_DFI_CLK_BUF;
    output [7:0] AXI_22_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_22_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_22_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_22_DFI_DW_RDDATA_VALID;
    output AXI_22_DFI_INIT_COMPLETE;
    output AXI_22_DFI_PHYUPD_REQ;
    output AXI_22_DFI_PHY_LP_STATE;
    output AXI_22_DFI_RST_N_BUF;
    output [5:0] AXI_22_MC_STATUS;
    output [7:0] AXI_22_PHY_STATUS;
    output [255:0] AXI_22_RDATA;
    output [31:0] AXI_22_RDATA_PARITY;
    output [5:0] AXI_22_RID;
    output AXI_22_RLAST;
    output [1:0] AXI_22_RRESP;
    output AXI_22_RVALID;
    output AXI_22_WREADY;
    output AXI_23_ARREADY;
    output AXI_23_AWREADY;
    output [5:0] AXI_23_BID;
    output [1:0] AXI_23_BRESP;
    output AXI_23_BVALID;
    output [1:0] AXI_23_DFI_AW_AERR_N;
    output AXI_23_DFI_CLK_BUF;
    output [7:0] AXI_23_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_23_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_23_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_23_DFI_DW_RDDATA_VALID;
    output AXI_23_DFI_INIT_COMPLETE;
    output AXI_23_DFI_PHYUPD_REQ;
    output AXI_23_DFI_PHY_LP_STATE;
    output AXI_23_DFI_RST_N_BUF;
    output [255:0] AXI_23_RDATA;
    output [31:0] AXI_23_RDATA_PARITY;
    output [5:0] AXI_23_RID;
    output AXI_23_RLAST;
    output [1:0] AXI_23_RRESP;
    output AXI_23_RVALID;
    output AXI_23_WREADY;
    output AXI_24_ARREADY;
    output AXI_24_AWREADY;
    output [5:0] AXI_24_BID;
    output [1:0] AXI_24_BRESP;
    output AXI_24_BVALID;
    output [1:0] AXI_24_DFI_AW_AERR_N;
    output AXI_24_DFI_CLK_BUF;
    output [7:0] AXI_24_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_24_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_24_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_24_DFI_DW_RDDATA_VALID;
    output AXI_24_DFI_INIT_COMPLETE;
    output AXI_24_DFI_PHYUPD_REQ;
    output AXI_24_DFI_PHY_LP_STATE;
    output AXI_24_DFI_RST_N_BUF;
    output [5:0] AXI_24_MC_STATUS;
    output [7:0] AXI_24_PHY_STATUS;
    output [255:0] AXI_24_RDATA;
    output [31:0] AXI_24_RDATA_PARITY;
    output [5:0] AXI_24_RID;
    output AXI_24_RLAST;
    output [1:0] AXI_24_RRESP;
    output AXI_24_RVALID;
    output AXI_24_WREADY;
    output AXI_25_ARREADY;
    output AXI_25_AWREADY;
    output [5:0] AXI_25_BID;
    output [1:0] AXI_25_BRESP;
    output AXI_25_BVALID;
    output [1:0] AXI_25_DFI_AW_AERR_N;
    output AXI_25_DFI_CLK_BUF;
    output [7:0] AXI_25_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_25_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_25_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_25_DFI_DW_RDDATA_VALID;
    output AXI_25_DFI_INIT_COMPLETE;
    output AXI_25_DFI_PHYUPD_REQ;
    output AXI_25_DFI_PHY_LP_STATE;
    output AXI_25_DFI_RST_N_BUF;
    output [255:0] AXI_25_RDATA;
    output [31:0] AXI_25_RDATA_PARITY;
    output [5:0] AXI_25_RID;
    output AXI_25_RLAST;
    output [1:0] AXI_25_RRESP;
    output AXI_25_RVALID;
    output AXI_25_WREADY;
    output AXI_26_ARREADY;
    output AXI_26_AWREADY;
    output [5:0] AXI_26_BID;
    output [1:0] AXI_26_BRESP;
    output AXI_26_BVALID;
    output [1:0] AXI_26_DFI_AW_AERR_N;
    output AXI_26_DFI_CLK_BUF;
    output [7:0] AXI_26_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_26_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_26_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_26_DFI_DW_RDDATA_VALID;
    output AXI_26_DFI_INIT_COMPLETE;
    output AXI_26_DFI_PHYUPD_REQ;
    output AXI_26_DFI_PHY_LP_STATE;
    output AXI_26_DFI_RST_N_BUF;
    output [5:0] AXI_26_MC_STATUS;
    output [7:0] AXI_26_PHY_STATUS;
    output [255:0] AXI_26_RDATA;
    output [31:0] AXI_26_RDATA_PARITY;
    output [5:0] AXI_26_RID;
    output AXI_26_RLAST;
    output [1:0] AXI_26_RRESP;
    output AXI_26_RVALID;
    output AXI_26_WREADY;
    output AXI_27_ARREADY;
    output AXI_27_AWREADY;
    output [5:0] AXI_27_BID;
    output [1:0] AXI_27_BRESP;
    output AXI_27_BVALID;
    output [1:0] AXI_27_DFI_AW_AERR_N;
    output AXI_27_DFI_CLK_BUF;
    output [7:0] AXI_27_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_27_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_27_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_27_DFI_DW_RDDATA_VALID;
    output AXI_27_DFI_INIT_COMPLETE;
    output AXI_27_DFI_PHYUPD_REQ;
    output AXI_27_DFI_PHY_LP_STATE;
    output AXI_27_DFI_RST_N_BUF;
    output [255:0] AXI_27_RDATA;
    output [31:0] AXI_27_RDATA_PARITY;
    output [5:0] AXI_27_RID;
    output AXI_27_RLAST;
    output [1:0] AXI_27_RRESP;
    output AXI_27_RVALID;
    output AXI_27_WREADY;
    output AXI_28_ARREADY;
    output AXI_28_AWREADY;
    output [5:0] AXI_28_BID;
    output [1:0] AXI_28_BRESP;
    output AXI_28_BVALID;
    output [1:0] AXI_28_DFI_AW_AERR_N;
    output AXI_28_DFI_CLK_BUF;
    output [7:0] AXI_28_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_28_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_28_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_28_DFI_DW_RDDATA_VALID;
    output AXI_28_DFI_INIT_COMPLETE;
    output AXI_28_DFI_PHYUPD_REQ;
    output AXI_28_DFI_PHY_LP_STATE;
    output AXI_28_DFI_RST_N_BUF;
    output [5:0] AXI_28_MC_STATUS;
    output [7:0] AXI_28_PHY_STATUS;
    output [255:0] AXI_28_RDATA;
    output [31:0] AXI_28_RDATA_PARITY;
    output [5:0] AXI_28_RID;
    output AXI_28_RLAST;
    output [1:0] AXI_28_RRESP;
    output AXI_28_RVALID;
    output AXI_28_WREADY;
    output AXI_29_ARREADY;
    output AXI_29_AWREADY;
    output [5:0] AXI_29_BID;
    output [1:0] AXI_29_BRESP;
    output AXI_29_BVALID;
    output [1:0] AXI_29_DFI_AW_AERR_N;
    output AXI_29_DFI_CLK_BUF;
    output [7:0] AXI_29_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_29_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_29_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_29_DFI_DW_RDDATA_VALID;
    output AXI_29_DFI_INIT_COMPLETE;
    output AXI_29_DFI_PHYUPD_REQ;
    output AXI_29_DFI_PHY_LP_STATE;
    output AXI_29_DFI_RST_N_BUF;
    output [255:0] AXI_29_RDATA;
    output [31:0] AXI_29_RDATA_PARITY;
    output [5:0] AXI_29_RID;
    output AXI_29_RLAST;
    output [1:0] AXI_29_RRESP;
    output AXI_29_RVALID;
    output AXI_29_WREADY;
    output AXI_30_ARREADY;
    output AXI_30_AWREADY;
    output [5:0] AXI_30_BID;
    output [1:0] AXI_30_BRESP;
    output AXI_30_BVALID;
    output [1:0] AXI_30_DFI_AW_AERR_N;
    output AXI_30_DFI_CLK_BUF;
    output [7:0] AXI_30_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_30_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_30_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_30_DFI_DW_RDDATA_VALID;
    output AXI_30_DFI_INIT_COMPLETE;
    output AXI_30_DFI_PHYUPD_REQ;
    output AXI_30_DFI_PHY_LP_STATE;
    output AXI_30_DFI_RST_N_BUF;
    output [5:0] AXI_30_MC_STATUS;
    output [7:0] AXI_30_PHY_STATUS;
    output [255:0] AXI_30_RDATA;
    output [31:0] AXI_30_RDATA_PARITY;
    output [5:0] AXI_30_RID;
    output AXI_30_RLAST;
    output [1:0] AXI_30_RRESP;
    output AXI_30_RVALID;
    output AXI_30_WREADY;
    output AXI_31_ARREADY;
    output AXI_31_AWREADY;
    output [5:0] AXI_31_BID;
    output [1:0] AXI_31_BRESP;
    output AXI_31_BVALID;
    output [1:0] AXI_31_DFI_AW_AERR_N;
    output AXI_31_DFI_CLK_BUF;
    output [7:0] AXI_31_DFI_DBI_BYTE_DISABLE;
    output [20:0] AXI_31_DFI_DW_RDDATA_DBI;
    output [7:0] AXI_31_DFI_DW_RDDATA_DERR;
    output [1:0] AXI_31_DFI_DW_RDDATA_VALID;
    output AXI_31_DFI_INIT_COMPLETE;
    output AXI_31_DFI_PHYUPD_REQ;
    output AXI_31_DFI_PHY_LP_STATE;
    output AXI_31_DFI_RST_N_BUF;
    output [255:0] AXI_31_RDATA;
    output [31:0] AXI_31_RDATA_PARITY;
    output [5:0] AXI_31_RID;
    output AXI_31_RLAST;
    output [1:0] AXI_31_RRESP;
    output AXI_31_RVALID;
    output AXI_31_WREADY;
    output DRAM_0_STAT_CATTRIP;
    output [2:0] DRAM_0_STAT_TEMP;
    output DRAM_1_STAT_CATTRIP;
    output [2:0] DRAM_1_STAT_TEMP;
    input [21:0] APB_0_PADDR;
    (* invertible_pin = "IS_APB_0_PCLK_INVERTED" *)
    input APB_0_PCLK;
    input APB_0_PENABLE;
    (* invertible_pin = "IS_APB_0_PRESET_N_INVERTED" *)
    input APB_0_PRESET_N;
    input APB_0_PSEL;
    input [31:0] APB_0_PWDATA;
    input APB_0_PWRITE;
    input [21:0] APB_1_PADDR;
    (* invertible_pin = "IS_APB_1_PCLK_INVERTED" *)
    input APB_1_PCLK;
    input APB_1_PENABLE;
    (* invertible_pin = "IS_APB_1_PRESET_N_INVERTED" *)
    input APB_1_PRESET_N;
    input APB_1_PSEL;
    input [31:0] APB_1_PWDATA;
    input APB_1_PWRITE;
    (* invertible_pin = "IS_AXI_00_ACLK_INVERTED" *)
    input AXI_00_ACLK;
    input [36:0] AXI_00_ARADDR;
    input [1:0] AXI_00_ARBURST;
    (* invertible_pin = "IS_AXI_00_ARESET_N_INVERTED" *)
    input AXI_00_ARESET_N;
    input [5:0] AXI_00_ARID;
    input [3:0] AXI_00_ARLEN;
    input [2:0] AXI_00_ARSIZE;
    input AXI_00_ARVALID;
    input [36:0] AXI_00_AWADDR;
    input [1:0] AXI_00_AWBURST;
    input [5:0] AXI_00_AWID;
    input [3:0] AXI_00_AWLEN;
    input [2:0] AXI_00_AWSIZE;
    input AXI_00_AWVALID;
    input AXI_00_BREADY;
    input AXI_00_DFI_LP_PWR_X_REQ;
    input AXI_00_RREADY;
    input [255:0] AXI_00_WDATA;
    input [31:0] AXI_00_WDATA_PARITY;
    input AXI_00_WLAST;
    input [31:0] AXI_00_WSTRB;
    input AXI_00_WVALID;
    (* invertible_pin = "IS_AXI_01_ACLK_INVERTED" *)
    input AXI_01_ACLK;
    input [36:0] AXI_01_ARADDR;
    input [1:0] AXI_01_ARBURST;
    (* invertible_pin = "IS_AXI_01_ARESET_N_INVERTED" *)
    input AXI_01_ARESET_N;
    input [5:0] AXI_01_ARID;
    input [3:0] AXI_01_ARLEN;
    input [2:0] AXI_01_ARSIZE;
    input AXI_01_ARVALID;
    input [36:0] AXI_01_AWADDR;
    input [1:0] AXI_01_AWBURST;
    input [5:0] AXI_01_AWID;
    input [3:0] AXI_01_AWLEN;
    input [2:0] AXI_01_AWSIZE;
    input AXI_01_AWVALID;
    input AXI_01_BREADY;
    input AXI_01_DFI_LP_PWR_X_REQ;
    input AXI_01_RREADY;
    input [255:0] AXI_01_WDATA;
    input [31:0] AXI_01_WDATA_PARITY;
    input AXI_01_WLAST;
    input [31:0] AXI_01_WSTRB;
    input AXI_01_WVALID;
    (* invertible_pin = "IS_AXI_02_ACLK_INVERTED" *)
    input AXI_02_ACLK;
    input [36:0] AXI_02_ARADDR;
    input [1:0] AXI_02_ARBURST;
    (* invertible_pin = "IS_AXI_02_ARESET_N_INVERTED" *)
    input AXI_02_ARESET_N;
    input [5:0] AXI_02_ARID;
    input [3:0] AXI_02_ARLEN;
    input [2:0] AXI_02_ARSIZE;
    input AXI_02_ARVALID;
    input [36:0] AXI_02_AWADDR;
    input [1:0] AXI_02_AWBURST;
    input [5:0] AXI_02_AWID;
    input [3:0] AXI_02_AWLEN;
    input [2:0] AXI_02_AWSIZE;
    input AXI_02_AWVALID;
    input AXI_02_BREADY;
    input AXI_02_DFI_LP_PWR_X_REQ;
    input AXI_02_RREADY;
    input [255:0] AXI_02_WDATA;
    input [31:0] AXI_02_WDATA_PARITY;
    input AXI_02_WLAST;
    input [31:0] AXI_02_WSTRB;
    input AXI_02_WVALID;
    (* invertible_pin = "IS_AXI_03_ACLK_INVERTED" *)
    input AXI_03_ACLK;
    input [36:0] AXI_03_ARADDR;
    input [1:0] AXI_03_ARBURST;
    (* invertible_pin = "IS_AXI_03_ARESET_N_INVERTED" *)
    input AXI_03_ARESET_N;
    input [5:0] AXI_03_ARID;
    input [3:0] AXI_03_ARLEN;
    input [2:0] AXI_03_ARSIZE;
    input AXI_03_ARVALID;
    input [36:0] AXI_03_AWADDR;
    input [1:0] AXI_03_AWBURST;
    input [5:0] AXI_03_AWID;
    input [3:0] AXI_03_AWLEN;
    input [2:0] AXI_03_AWSIZE;
    input AXI_03_AWVALID;
    input AXI_03_BREADY;
    input AXI_03_DFI_LP_PWR_X_REQ;
    input AXI_03_RREADY;
    input [255:0] AXI_03_WDATA;
    input [31:0] AXI_03_WDATA_PARITY;
    input AXI_03_WLAST;
    input [31:0] AXI_03_WSTRB;
    input AXI_03_WVALID;
    (* invertible_pin = "IS_AXI_04_ACLK_INVERTED" *)
    input AXI_04_ACLK;
    input [36:0] AXI_04_ARADDR;
    input [1:0] AXI_04_ARBURST;
    (* invertible_pin = "IS_AXI_04_ARESET_N_INVERTED" *)
    input AXI_04_ARESET_N;
    input [5:0] AXI_04_ARID;
    input [3:0] AXI_04_ARLEN;
    input [2:0] AXI_04_ARSIZE;
    input AXI_04_ARVALID;
    input [36:0] AXI_04_AWADDR;
    input [1:0] AXI_04_AWBURST;
    input [5:0] AXI_04_AWID;
    input [3:0] AXI_04_AWLEN;
    input [2:0] AXI_04_AWSIZE;
    input AXI_04_AWVALID;
    input AXI_04_BREADY;
    input AXI_04_DFI_LP_PWR_X_REQ;
    input AXI_04_RREADY;
    input [255:0] AXI_04_WDATA;
    input [31:0] AXI_04_WDATA_PARITY;
    input AXI_04_WLAST;
    input [31:0] AXI_04_WSTRB;
    input AXI_04_WVALID;
    (* invertible_pin = "IS_AXI_05_ACLK_INVERTED" *)
    input AXI_05_ACLK;
    input [36:0] AXI_05_ARADDR;
    input [1:0] AXI_05_ARBURST;
    (* invertible_pin = "IS_AXI_05_ARESET_N_INVERTED" *)
    input AXI_05_ARESET_N;
    input [5:0] AXI_05_ARID;
    input [3:0] AXI_05_ARLEN;
    input [2:0] AXI_05_ARSIZE;
    input AXI_05_ARVALID;
    input [36:0] AXI_05_AWADDR;
    input [1:0] AXI_05_AWBURST;
    input [5:0] AXI_05_AWID;
    input [3:0] AXI_05_AWLEN;
    input [2:0] AXI_05_AWSIZE;
    input AXI_05_AWVALID;
    input AXI_05_BREADY;
    input AXI_05_DFI_LP_PWR_X_REQ;
    input AXI_05_RREADY;
    input [255:0] AXI_05_WDATA;
    input [31:0] AXI_05_WDATA_PARITY;
    input AXI_05_WLAST;
    input [31:0] AXI_05_WSTRB;
    input AXI_05_WVALID;
    (* invertible_pin = "IS_AXI_06_ACLK_INVERTED" *)
    input AXI_06_ACLK;
    input [36:0] AXI_06_ARADDR;
    input [1:0] AXI_06_ARBURST;
    (* invertible_pin = "IS_AXI_06_ARESET_N_INVERTED" *)
    input AXI_06_ARESET_N;
    input [5:0] AXI_06_ARID;
    input [3:0] AXI_06_ARLEN;
    input [2:0] AXI_06_ARSIZE;
    input AXI_06_ARVALID;
    input [36:0] AXI_06_AWADDR;
    input [1:0] AXI_06_AWBURST;
    input [5:0] AXI_06_AWID;
    input [3:0] AXI_06_AWLEN;
    input [2:0] AXI_06_AWSIZE;
    input AXI_06_AWVALID;
    input AXI_06_BREADY;
    input AXI_06_DFI_LP_PWR_X_REQ;
    input AXI_06_RREADY;
    input [255:0] AXI_06_WDATA;
    input [31:0] AXI_06_WDATA_PARITY;
    input AXI_06_WLAST;
    input [31:0] AXI_06_WSTRB;
    input AXI_06_WVALID;
    (* invertible_pin = "IS_AXI_07_ACLK_INVERTED" *)
    input AXI_07_ACLK;
    input [36:0] AXI_07_ARADDR;
    input [1:0] AXI_07_ARBURST;
    (* invertible_pin = "IS_AXI_07_ARESET_N_INVERTED" *)
    input AXI_07_ARESET_N;
    input [5:0] AXI_07_ARID;
    input [3:0] AXI_07_ARLEN;
    input [2:0] AXI_07_ARSIZE;
    input AXI_07_ARVALID;
    input [36:0] AXI_07_AWADDR;
    input [1:0] AXI_07_AWBURST;
    input [5:0] AXI_07_AWID;
    input [3:0] AXI_07_AWLEN;
    input [2:0] AXI_07_AWSIZE;
    input AXI_07_AWVALID;
    input AXI_07_BREADY;
    input AXI_07_DFI_LP_PWR_X_REQ;
    input AXI_07_RREADY;
    input [255:0] AXI_07_WDATA;
    input [31:0] AXI_07_WDATA_PARITY;
    input AXI_07_WLAST;
    input [31:0] AXI_07_WSTRB;
    input AXI_07_WVALID;
    (* invertible_pin = "IS_AXI_08_ACLK_INVERTED" *)
    input AXI_08_ACLK;
    input [36:0] AXI_08_ARADDR;
    input [1:0] AXI_08_ARBURST;
    (* invertible_pin = "IS_AXI_08_ARESET_N_INVERTED" *)
    input AXI_08_ARESET_N;
    input [5:0] AXI_08_ARID;
    input [3:0] AXI_08_ARLEN;
    input [2:0] AXI_08_ARSIZE;
    input AXI_08_ARVALID;
    input [36:0] AXI_08_AWADDR;
    input [1:0] AXI_08_AWBURST;
    input [5:0] AXI_08_AWID;
    input [3:0] AXI_08_AWLEN;
    input [2:0] AXI_08_AWSIZE;
    input AXI_08_AWVALID;
    input AXI_08_BREADY;
    input AXI_08_DFI_LP_PWR_X_REQ;
    input AXI_08_RREADY;
    input [255:0] AXI_08_WDATA;
    input [31:0] AXI_08_WDATA_PARITY;
    input AXI_08_WLAST;
    input [31:0] AXI_08_WSTRB;
    input AXI_08_WVALID;
    (* invertible_pin = "IS_AXI_09_ACLK_INVERTED" *)
    input AXI_09_ACLK;
    input [36:0] AXI_09_ARADDR;
    input [1:0] AXI_09_ARBURST;
    (* invertible_pin = "IS_AXI_09_ARESET_N_INVERTED" *)
    input AXI_09_ARESET_N;
    input [5:0] AXI_09_ARID;
    input [3:0] AXI_09_ARLEN;
    input [2:0] AXI_09_ARSIZE;
    input AXI_09_ARVALID;
    input [36:0] AXI_09_AWADDR;
    input [1:0] AXI_09_AWBURST;
    input [5:0] AXI_09_AWID;
    input [3:0] AXI_09_AWLEN;
    input [2:0] AXI_09_AWSIZE;
    input AXI_09_AWVALID;
    input AXI_09_BREADY;
    input AXI_09_DFI_LP_PWR_X_REQ;
    input AXI_09_RREADY;
    input [255:0] AXI_09_WDATA;
    input [31:0] AXI_09_WDATA_PARITY;
    input AXI_09_WLAST;
    input [31:0] AXI_09_WSTRB;
    input AXI_09_WVALID;
    (* invertible_pin = "IS_AXI_10_ACLK_INVERTED" *)
    input AXI_10_ACLK;
    input [36:0] AXI_10_ARADDR;
    input [1:0] AXI_10_ARBURST;
    (* invertible_pin = "IS_AXI_10_ARESET_N_INVERTED" *)
    input AXI_10_ARESET_N;
    input [5:0] AXI_10_ARID;
    input [3:0] AXI_10_ARLEN;
    input [2:0] AXI_10_ARSIZE;
    input AXI_10_ARVALID;
    input [36:0] AXI_10_AWADDR;
    input [1:0] AXI_10_AWBURST;
    input [5:0] AXI_10_AWID;
    input [3:0] AXI_10_AWLEN;
    input [2:0] AXI_10_AWSIZE;
    input AXI_10_AWVALID;
    input AXI_10_BREADY;
    input AXI_10_DFI_LP_PWR_X_REQ;
    input AXI_10_RREADY;
    input [255:0] AXI_10_WDATA;
    input [31:0] AXI_10_WDATA_PARITY;
    input AXI_10_WLAST;
    input [31:0] AXI_10_WSTRB;
    input AXI_10_WVALID;
    (* invertible_pin = "IS_AXI_11_ACLK_INVERTED" *)
    input AXI_11_ACLK;
    input [36:0] AXI_11_ARADDR;
    input [1:0] AXI_11_ARBURST;
    (* invertible_pin = "IS_AXI_11_ARESET_N_INVERTED" *)
    input AXI_11_ARESET_N;
    input [5:0] AXI_11_ARID;
    input [3:0] AXI_11_ARLEN;
    input [2:0] AXI_11_ARSIZE;
    input AXI_11_ARVALID;
    input [36:0] AXI_11_AWADDR;
    input [1:0] AXI_11_AWBURST;
    input [5:0] AXI_11_AWID;
    input [3:0] AXI_11_AWLEN;
    input [2:0] AXI_11_AWSIZE;
    input AXI_11_AWVALID;
    input AXI_11_BREADY;
    input AXI_11_DFI_LP_PWR_X_REQ;
    input AXI_11_RREADY;
    input [255:0] AXI_11_WDATA;
    input [31:0] AXI_11_WDATA_PARITY;
    input AXI_11_WLAST;
    input [31:0] AXI_11_WSTRB;
    input AXI_11_WVALID;
    (* invertible_pin = "IS_AXI_12_ACLK_INVERTED" *)
    input AXI_12_ACLK;
    input [36:0] AXI_12_ARADDR;
    input [1:0] AXI_12_ARBURST;
    (* invertible_pin = "IS_AXI_12_ARESET_N_INVERTED" *)
    input AXI_12_ARESET_N;
    input [5:0] AXI_12_ARID;
    input [3:0] AXI_12_ARLEN;
    input [2:0] AXI_12_ARSIZE;
    input AXI_12_ARVALID;
    input [36:0] AXI_12_AWADDR;
    input [1:0] AXI_12_AWBURST;
    input [5:0] AXI_12_AWID;
    input [3:0] AXI_12_AWLEN;
    input [2:0] AXI_12_AWSIZE;
    input AXI_12_AWVALID;
    input AXI_12_BREADY;
    input AXI_12_DFI_LP_PWR_X_REQ;
    input AXI_12_RREADY;
    input [255:0] AXI_12_WDATA;
    input [31:0] AXI_12_WDATA_PARITY;
    input AXI_12_WLAST;
    input [31:0] AXI_12_WSTRB;
    input AXI_12_WVALID;
    (* invertible_pin = "IS_AXI_13_ACLK_INVERTED" *)
    input AXI_13_ACLK;
    input [36:0] AXI_13_ARADDR;
    input [1:0] AXI_13_ARBURST;
    (* invertible_pin = "IS_AXI_13_ARESET_N_INVERTED" *)
    input AXI_13_ARESET_N;
    input [5:0] AXI_13_ARID;
    input [3:0] AXI_13_ARLEN;
    input [2:0] AXI_13_ARSIZE;
    input AXI_13_ARVALID;
    input [36:0] AXI_13_AWADDR;
    input [1:0] AXI_13_AWBURST;
    input [5:0] AXI_13_AWID;
    input [3:0] AXI_13_AWLEN;
    input [2:0] AXI_13_AWSIZE;
    input AXI_13_AWVALID;
    input AXI_13_BREADY;
    input AXI_13_DFI_LP_PWR_X_REQ;
    input AXI_13_RREADY;
    input [255:0] AXI_13_WDATA;
    input [31:0] AXI_13_WDATA_PARITY;
    input AXI_13_WLAST;
    input [31:0] AXI_13_WSTRB;
    input AXI_13_WVALID;
    (* invertible_pin = "IS_AXI_14_ACLK_INVERTED" *)
    input AXI_14_ACLK;
    input [36:0] AXI_14_ARADDR;
    input [1:0] AXI_14_ARBURST;
    (* invertible_pin = "IS_AXI_14_ARESET_N_INVERTED" *)
    input AXI_14_ARESET_N;
    input [5:0] AXI_14_ARID;
    input [3:0] AXI_14_ARLEN;
    input [2:0] AXI_14_ARSIZE;
    input AXI_14_ARVALID;
    input [36:0] AXI_14_AWADDR;
    input [1:0] AXI_14_AWBURST;
    input [5:0] AXI_14_AWID;
    input [3:0] AXI_14_AWLEN;
    input [2:0] AXI_14_AWSIZE;
    input AXI_14_AWVALID;
    input AXI_14_BREADY;
    input AXI_14_DFI_LP_PWR_X_REQ;
    input AXI_14_RREADY;
    input [255:0] AXI_14_WDATA;
    input [31:0] AXI_14_WDATA_PARITY;
    input AXI_14_WLAST;
    input [31:0] AXI_14_WSTRB;
    input AXI_14_WVALID;
    (* invertible_pin = "IS_AXI_15_ACLK_INVERTED" *)
    input AXI_15_ACLK;
    input [36:0] AXI_15_ARADDR;
    input [1:0] AXI_15_ARBURST;
    (* invertible_pin = "IS_AXI_15_ARESET_N_INVERTED" *)
    input AXI_15_ARESET_N;
    input [5:0] AXI_15_ARID;
    input [3:0] AXI_15_ARLEN;
    input [2:0] AXI_15_ARSIZE;
    input AXI_15_ARVALID;
    input [36:0] AXI_15_AWADDR;
    input [1:0] AXI_15_AWBURST;
    input [5:0] AXI_15_AWID;
    input [3:0] AXI_15_AWLEN;
    input [2:0] AXI_15_AWSIZE;
    input AXI_15_AWVALID;
    input AXI_15_BREADY;
    input AXI_15_DFI_LP_PWR_X_REQ;
    input AXI_15_RREADY;
    input [255:0] AXI_15_WDATA;
    input [31:0] AXI_15_WDATA_PARITY;
    input AXI_15_WLAST;
    input [31:0] AXI_15_WSTRB;
    input AXI_15_WVALID;
    (* invertible_pin = "IS_AXI_16_ACLK_INVERTED" *)
    input AXI_16_ACLK;
    input [36:0] AXI_16_ARADDR;
    input [1:0] AXI_16_ARBURST;
    (* invertible_pin = "IS_AXI_16_ARESET_N_INVERTED" *)
    input AXI_16_ARESET_N;
    input [5:0] AXI_16_ARID;
    input [3:0] AXI_16_ARLEN;
    input [2:0] AXI_16_ARSIZE;
    input AXI_16_ARVALID;
    input [36:0] AXI_16_AWADDR;
    input [1:0] AXI_16_AWBURST;
    input [5:0] AXI_16_AWID;
    input [3:0] AXI_16_AWLEN;
    input [2:0] AXI_16_AWSIZE;
    input AXI_16_AWVALID;
    input AXI_16_BREADY;
    input AXI_16_DFI_LP_PWR_X_REQ;
    input AXI_16_RREADY;
    input [255:0] AXI_16_WDATA;
    input [31:0] AXI_16_WDATA_PARITY;
    input AXI_16_WLAST;
    input [31:0] AXI_16_WSTRB;
    input AXI_16_WVALID;
    (* invertible_pin = "IS_AXI_17_ACLK_INVERTED" *)
    input AXI_17_ACLK;
    input [36:0] AXI_17_ARADDR;
    input [1:0] AXI_17_ARBURST;
    (* invertible_pin = "IS_AXI_17_ARESET_N_INVERTED" *)
    input AXI_17_ARESET_N;
    input [5:0] AXI_17_ARID;
    input [3:0] AXI_17_ARLEN;
    input [2:0] AXI_17_ARSIZE;
    input AXI_17_ARVALID;
    input [36:0] AXI_17_AWADDR;
    input [1:0] AXI_17_AWBURST;
    input [5:0] AXI_17_AWID;
    input [3:0] AXI_17_AWLEN;
    input [2:0] AXI_17_AWSIZE;
    input AXI_17_AWVALID;
    input AXI_17_BREADY;
    input AXI_17_DFI_LP_PWR_X_REQ;
    input AXI_17_RREADY;
    input [255:0] AXI_17_WDATA;
    input [31:0] AXI_17_WDATA_PARITY;
    input AXI_17_WLAST;
    input [31:0] AXI_17_WSTRB;
    input AXI_17_WVALID;
    (* invertible_pin = "IS_AXI_18_ACLK_INVERTED" *)
    input AXI_18_ACLK;
    input [36:0] AXI_18_ARADDR;
    input [1:0] AXI_18_ARBURST;
    (* invertible_pin = "IS_AXI_18_ARESET_N_INVERTED" *)
    input AXI_18_ARESET_N;
    input [5:0] AXI_18_ARID;
    input [3:0] AXI_18_ARLEN;
    input [2:0] AXI_18_ARSIZE;
    input AXI_18_ARVALID;
    input [36:0] AXI_18_AWADDR;
    input [1:0] AXI_18_AWBURST;
    input [5:0] AXI_18_AWID;
    input [3:0] AXI_18_AWLEN;
    input [2:0] AXI_18_AWSIZE;
    input AXI_18_AWVALID;
    input AXI_18_BREADY;
    input AXI_18_DFI_LP_PWR_X_REQ;
    input AXI_18_RREADY;
    input [255:0] AXI_18_WDATA;
    input [31:0] AXI_18_WDATA_PARITY;
    input AXI_18_WLAST;
    input [31:0] AXI_18_WSTRB;
    input AXI_18_WVALID;
    (* invertible_pin = "IS_AXI_19_ACLK_INVERTED" *)
    input AXI_19_ACLK;
    input [36:0] AXI_19_ARADDR;
    input [1:0] AXI_19_ARBURST;
    (* invertible_pin = "IS_AXI_19_ARESET_N_INVERTED" *)
    input AXI_19_ARESET_N;
    input [5:0] AXI_19_ARID;
    input [3:0] AXI_19_ARLEN;
    input [2:0] AXI_19_ARSIZE;
    input AXI_19_ARVALID;
    input [36:0] AXI_19_AWADDR;
    input [1:0] AXI_19_AWBURST;
    input [5:0] AXI_19_AWID;
    input [3:0] AXI_19_AWLEN;
    input [2:0] AXI_19_AWSIZE;
    input AXI_19_AWVALID;
    input AXI_19_BREADY;
    input AXI_19_DFI_LP_PWR_X_REQ;
    input AXI_19_RREADY;
    input [255:0] AXI_19_WDATA;
    input [31:0] AXI_19_WDATA_PARITY;
    input AXI_19_WLAST;
    input [31:0] AXI_19_WSTRB;
    input AXI_19_WVALID;
    (* invertible_pin = "IS_AXI_20_ACLK_INVERTED" *)
    input AXI_20_ACLK;
    input [36:0] AXI_20_ARADDR;
    input [1:0] AXI_20_ARBURST;
    (* invertible_pin = "IS_AXI_20_ARESET_N_INVERTED" *)
    input AXI_20_ARESET_N;
    input [5:0] AXI_20_ARID;
    input [3:0] AXI_20_ARLEN;
    input [2:0] AXI_20_ARSIZE;
    input AXI_20_ARVALID;
    input [36:0] AXI_20_AWADDR;
    input [1:0] AXI_20_AWBURST;
    input [5:0] AXI_20_AWID;
    input [3:0] AXI_20_AWLEN;
    input [2:0] AXI_20_AWSIZE;
    input AXI_20_AWVALID;
    input AXI_20_BREADY;
    input AXI_20_DFI_LP_PWR_X_REQ;
    input AXI_20_RREADY;
    input [255:0] AXI_20_WDATA;
    input [31:0] AXI_20_WDATA_PARITY;
    input AXI_20_WLAST;
    input [31:0] AXI_20_WSTRB;
    input AXI_20_WVALID;
    (* invertible_pin = "IS_AXI_21_ACLK_INVERTED" *)
    input AXI_21_ACLK;
    input [36:0] AXI_21_ARADDR;
    input [1:0] AXI_21_ARBURST;
    (* invertible_pin = "IS_AXI_21_ARESET_N_INVERTED" *)
    input AXI_21_ARESET_N;
    input [5:0] AXI_21_ARID;
    input [3:0] AXI_21_ARLEN;
    input [2:0] AXI_21_ARSIZE;
    input AXI_21_ARVALID;
    input [36:0] AXI_21_AWADDR;
    input [1:0] AXI_21_AWBURST;
    input [5:0] AXI_21_AWID;
    input [3:0] AXI_21_AWLEN;
    input [2:0] AXI_21_AWSIZE;
    input AXI_21_AWVALID;
    input AXI_21_BREADY;
    input AXI_21_DFI_LP_PWR_X_REQ;
    input AXI_21_RREADY;
    input [255:0] AXI_21_WDATA;
    input [31:0] AXI_21_WDATA_PARITY;
    input AXI_21_WLAST;
    input [31:0] AXI_21_WSTRB;
    input AXI_21_WVALID;
    (* invertible_pin = "IS_AXI_22_ACLK_INVERTED" *)
    input AXI_22_ACLK;
    input [36:0] AXI_22_ARADDR;
    input [1:0] AXI_22_ARBURST;
    (* invertible_pin = "IS_AXI_22_ARESET_N_INVERTED" *)
    input AXI_22_ARESET_N;
    input [5:0] AXI_22_ARID;
    input [3:0] AXI_22_ARLEN;
    input [2:0] AXI_22_ARSIZE;
    input AXI_22_ARVALID;
    input [36:0] AXI_22_AWADDR;
    input [1:0] AXI_22_AWBURST;
    input [5:0] AXI_22_AWID;
    input [3:0] AXI_22_AWLEN;
    input [2:0] AXI_22_AWSIZE;
    input AXI_22_AWVALID;
    input AXI_22_BREADY;
    input AXI_22_DFI_LP_PWR_X_REQ;
    input AXI_22_RREADY;
    input [255:0] AXI_22_WDATA;
    input [31:0] AXI_22_WDATA_PARITY;
    input AXI_22_WLAST;
    input [31:0] AXI_22_WSTRB;
    input AXI_22_WVALID;
    (* invertible_pin = "IS_AXI_23_ACLK_INVERTED" *)
    input AXI_23_ACLK;
    input [36:0] AXI_23_ARADDR;
    input [1:0] AXI_23_ARBURST;
    (* invertible_pin = "IS_AXI_23_ARESET_N_INVERTED" *)
    input AXI_23_ARESET_N;
    input [5:0] AXI_23_ARID;
    input [3:0] AXI_23_ARLEN;
    input [2:0] AXI_23_ARSIZE;
    input AXI_23_ARVALID;
    input [36:0] AXI_23_AWADDR;
    input [1:0] AXI_23_AWBURST;
    input [5:0] AXI_23_AWID;
    input [3:0] AXI_23_AWLEN;
    input [2:0] AXI_23_AWSIZE;
    input AXI_23_AWVALID;
    input AXI_23_BREADY;
    input AXI_23_DFI_LP_PWR_X_REQ;
    input AXI_23_RREADY;
    input [255:0] AXI_23_WDATA;
    input [31:0] AXI_23_WDATA_PARITY;
    input AXI_23_WLAST;
    input [31:0] AXI_23_WSTRB;
    input AXI_23_WVALID;
    (* invertible_pin = "IS_AXI_24_ACLK_INVERTED" *)
    input AXI_24_ACLK;
    input [36:0] AXI_24_ARADDR;
    input [1:0] AXI_24_ARBURST;
    (* invertible_pin = "IS_AXI_24_ARESET_N_INVERTED" *)
    input AXI_24_ARESET_N;
    input [5:0] AXI_24_ARID;
    input [3:0] AXI_24_ARLEN;
    input [2:0] AXI_24_ARSIZE;
    input AXI_24_ARVALID;
    input [36:0] AXI_24_AWADDR;
    input [1:0] AXI_24_AWBURST;
    input [5:0] AXI_24_AWID;
    input [3:0] AXI_24_AWLEN;
    input [2:0] AXI_24_AWSIZE;
    input AXI_24_AWVALID;
    input AXI_24_BREADY;
    input AXI_24_DFI_LP_PWR_X_REQ;
    input AXI_24_RREADY;
    input [255:0] AXI_24_WDATA;
    input [31:0] AXI_24_WDATA_PARITY;
    input AXI_24_WLAST;
    input [31:0] AXI_24_WSTRB;
    input AXI_24_WVALID;
    (* invertible_pin = "IS_AXI_25_ACLK_INVERTED" *)
    input AXI_25_ACLK;
    input [36:0] AXI_25_ARADDR;
    input [1:0] AXI_25_ARBURST;
    (* invertible_pin = "IS_AXI_25_ARESET_N_INVERTED" *)
    input AXI_25_ARESET_N;
    input [5:0] AXI_25_ARID;
    input [3:0] AXI_25_ARLEN;
    input [2:0] AXI_25_ARSIZE;
    input AXI_25_ARVALID;
    input [36:0] AXI_25_AWADDR;
    input [1:0] AXI_25_AWBURST;
    input [5:0] AXI_25_AWID;
    input [3:0] AXI_25_AWLEN;
    input [2:0] AXI_25_AWSIZE;
    input AXI_25_AWVALID;
    input AXI_25_BREADY;
    input AXI_25_DFI_LP_PWR_X_REQ;
    input AXI_25_RREADY;
    input [255:0] AXI_25_WDATA;
    input [31:0] AXI_25_WDATA_PARITY;
    input AXI_25_WLAST;
    input [31:0] AXI_25_WSTRB;
    input AXI_25_WVALID;
    (* invertible_pin = "IS_AXI_26_ACLK_INVERTED" *)
    input AXI_26_ACLK;
    input [36:0] AXI_26_ARADDR;
    input [1:0] AXI_26_ARBURST;
    (* invertible_pin = "IS_AXI_26_ARESET_N_INVERTED" *)
    input AXI_26_ARESET_N;
    input [5:0] AXI_26_ARID;
    input [3:0] AXI_26_ARLEN;
    input [2:0] AXI_26_ARSIZE;
    input AXI_26_ARVALID;
    input [36:0] AXI_26_AWADDR;
    input [1:0] AXI_26_AWBURST;
    input [5:0] AXI_26_AWID;
    input [3:0] AXI_26_AWLEN;
    input [2:0] AXI_26_AWSIZE;
    input AXI_26_AWVALID;
    input AXI_26_BREADY;
    input AXI_26_DFI_LP_PWR_X_REQ;
    input AXI_26_RREADY;
    input [255:0] AXI_26_WDATA;
    input [31:0] AXI_26_WDATA_PARITY;
    input AXI_26_WLAST;
    input [31:0] AXI_26_WSTRB;
    input AXI_26_WVALID;
    (* invertible_pin = "IS_AXI_27_ACLK_INVERTED" *)
    input AXI_27_ACLK;
    input [36:0] AXI_27_ARADDR;
    input [1:0] AXI_27_ARBURST;
    (* invertible_pin = "IS_AXI_27_ARESET_N_INVERTED" *)
    input AXI_27_ARESET_N;
    input [5:0] AXI_27_ARID;
    input [3:0] AXI_27_ARLEN;
    input [2:0] AXI_27_ARSIZE;
    input AXI_27_ARVALID;
    input [36:0] AXI_27_AWADDR;
    input [1:0] AXI_27_AWBURST;
    input [5:0] AXI_27_AWID;
    input [3:0] AXI_27_AWLEN;
    input [2:0] AXI_27_AWSIZE;
    input AXI_27_AWVALID;
    input AXI_27_BREADY;
    input AXI_27_DFI_LP_PWR_X_REQ;
    input AXI_27_RREADY;
    input [255:0] AXI_27_WDATA;
    input [31:0] AXI_27_WDATA_PARITY;
    input AXI_27_WLAST;
    input [31:0] AXI_27_WSTRB;
    input AXI_27_WVALID;
    (* invertible_pin = "IS_AXI_28_ACLK_INVERTED" *)
    input AXI_28_ACLK;
    input [36:0] AXI_28_ARADDR;
    input [1:0] AXI_28_ARBURST;
    (* invertible_pin = "IS_AXI_28_ARESET_N_INVERTED" *)
    input AXI_28_ARESET_N;
    input [5:0] AXI_28_ARID;
    input [3:0] AXI_28_ARLEN;
    input [2:0] AXI_28_ARSIZE;
    input AXI_28_ARVALID;
    input [36:0] AXI_28_AWADDR;
    input [1:0] AXI_28_AWBURST;
    input [5:0] AXI_28_AWID;
    input [3:0] AXI_28_AWLEN;
    input [2:0] AXI_28_AWSIZE;
    input AXI_28_AWVALID;
    input AXI_28_BREADY;
    input AXI_28_DFI_LP_PWR_X_REQ;
    input AXI_28_RREADY;
    input [255:0] AXI_28_WDATA;
    input [31:0] AXI_28_WDATA_PARITY;
    input AXI_28_WLAST;
    input [31:0] AXI_28_WSTRB;
    input AXI_28_WVALID;
    (* invertible_pin = "IS_AXI_29_ACLK_INVERTED" *)
    input AXI_29_ACLK;
    input [36:0] AXI_29_ARADDR;
    input [1:0] AXI_29_ARBURST;
    (* invertible_pin = "IS_AXI_29_ARESET_N_INVERTED" *)
    input AXI_29_ARESET_N;
    input [5:0] AXI_29_ARID;
    input [3:0] AXI_29_ARLEN;
    input [2:0] AXI_29_ARSIZE;
    input AXI_29_ARVALID;
    input [36:0] AXI_29_AWADDR;
    input [1:0] AXI_29_AWBURST;
    input [5:0] AXI_29_AWID;
    input [3:0] AXI_29_AWLEN;
    input [2:0] AXI_29_AWSIZE;
    input AXI_29_AWVALID;
    input AXI_29_BREADY;
    input AXI_29_DFI_LP_PWR_X_REQ;
    input AXI_29_RREADY;
    input [255:0] AXI_29_WDATA;
    input [31:0] AXI_29_WDATA_PARITY;
    input AXI_29_WLAST;
    input [31:0] AXI_29_WSTRB;
    input AXI_29_WVALID;
    (* invertible_pin = "IS_AXI_30_ACLK_INVERTED" *)
    input AXI_30_ACLK;
    input [36:0] AXI_30_ARADDR;
    input [1:0] AXI_30_ARBURST;
    (* invertible_pin = "IS_AXI_30_ARESET_N_INVERTED" *)
    input AXI_30_ARESET_N;
    input [5:0] AXI_30_ARID;
    input [3:0] AXI_30_ARLEN;
    input [2:0] AXI_30_ARSIZE;
    input AXI_30_ARVALID;
    input [36:0] AXI_30_AWADDR;
    input [1:0] AXI_30_AWBURST;
    input [5:0] AXI_30_AWID;
    input [3:0] AXI_30_AWLEN;
    input [2:0] AXI_30_AWSIZE;
    input AXI_30_AWVALID;
    input AXI_30_BREADY;
    input AXI_30_DFI_LP_PWR_X_REQ;
    input AXI_30_RREADY;
    input [255:0] AXI_30_WDATA;
    input [31:0] AXI_30_WDATA_PARITY;
    input AXI_30_WLAST;
    input [31:0] AXI_30_WSTRB;
    input AXI_30_WVALID;
    (* invertible_pin = "IS_AXI_31_ACLK_INVERTED" *)
    input AXI_31_ACLK;
    input [36:0] AXI_31_ARADDR;
    input [1:0] AXI_31_ARBURST;
    (* invertible_pin = "IS_AXI_31_ARESET_N_INVERTED" *)
    input AXI_31_ARESET_N;
    input [5:0] AXI_31_ARID;
    input [3:0] AXI_31_ARLEN;
    input [2:0] AXI_31_ARSIZE;
    input AXI_31_ARVALID;
    input [36:0] AXI_31_AWADDR;
    input [1:0] AXI_31_AWBURST;
    input [5:0] AXI_31_AWID;
    input [3:0] AXI_31_AWLEN;
    input [2:0] AXI_31_AWSIZE;
    input AXI_31_AWVALID;
    input AXI_31_BREADY;
    input AXI_31_DFI_LP_PWR_X_REQ;
    input AXI_31_RREADY;
    input [255:0] AXI_31_WDATA;
    input [31:0] AXI_31_WDATA_PARITY;
    input AXI_31_WLAST;
    input [31:0] AXI_31_WSTRB;
    input AXI_31_WVALID;
    input BSCAN_DRCK_0;
    input BSCAN_DRCK_1;
    input BSCAN_TCK_0;
    input BSCAN_TCK_1;
    input HBM_REF_CLK_0;
    input HBM_REF_CLK_1;
    input MBIST_EN_00;
    input MBIST_EN_01;
    input MBIST_EN_02;
    input MBIST_EN_03;
    input MBIST_EN_04;
    input MBIST_EN_05;
    input MBIST_EN_06;
    input MBIST_EN_07;
    input MBIST_EN_08;
    input MBIST_EN_09;
    input MBIST_EN_10;
    input MBIST_EN_11;
    input MBIST_EN_12;
    input MBIST_EN_13;
    input MBIST_EN_14;
    input MBIST_EN_15;
endmodule

module ILKN (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "TRUE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0000;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0008;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "TRUE";
    parameter [6:0] CTL_TX_FC_CALLEN = 7'h00;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_VERSION = "2.0";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

module ILKNE4 (...);
    parameter BYPASS = "FALSE";
    parameter [1:0] CTL_RX_BURSTMAX = 2'h3;
    parameter [1:0] CTL_RX_CHAN_EXT = 2'h0;
    parameter [3:0] CTL_RX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_RX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter CTL_RX_PACKET_MODE = "FALSE";
    parameter [2:0] CTL_RX_RETRANS_MULT = 3'h0;
    parameter [3:0] CTL_RX_RETRANS_RETRY = 4'h2;
    parameter [15:0] CTL_RX_RETRANS_TIMER1 = 16'h0009;
    parameter [15:0] CTL_RX_RETRANS_TIMER2 = 16'h0000;
    parameter [11:0] CTL_RX_RETRANS_WDOG = 12'h000;
    parameter [7:0] CTL_RX_RETRANS_WRAP_TIMER = 8'h00;
    parameter CTL_TEST_MODE_PIN_CHAR = "FALSE";
    parameter [1:0] CTL_TX_BURSTMAX = 2'h3;
    parameter [2:0] CTL_TX_BURSTSHORT = 3'h1;
    parameter [1:0] CTL_TX_CHAN_EXT = 2'h0;
    parameter CTL_TX_DISABLE_SKIPWORD = "FALSE";
    parameter [3:0] CTL_TX_FC_CALLEN = 4'hF;
    parameter [3:0] CTL_TX_LAST_LANE = 4'hB;
    parameter [15:0] CTL_TX_MFRAMELEN_MINUS1 = 16'h07FF;
    parameter [13:0] CTL_TX_RETRANS_DEPTH = 14'h0800;
    parameter [2:0] CTL_TX_RETRANS_MULT = 3'h0;
    parameter [1:0] CTL_TX_RETRANS_RAM_BANKS = 2'h3;
    parameter MODE = "TRUE";
    parameter SIM_DEVICE = "ULTRASCALE_PLUS";
    parameter TEST_MODE_PIN_CHAR = "FALSE";
    output [15:0] DRP_DO;
    output DRP_RDY;
    output [65:0] RX_BYPASS_DATAOUT00;
    output [65:0] RX_BYPASS_DATAOUT01;
    output [65:0] RX_BYPASS_DATAOUT02;
    output [65:0] RX_BYPASS_DATAOUT03;
    output [65:0] RX_BYPASS_DATAOUT04;
    output [65:0] RX_BYPASS_DATAOUT05;
    output [65:0] RX_BYPASS_DATAOUT06;
    output [65:0] RX_BYPASS_DATAOUT07;
    output [65:0] RX_BYPASS_DATAOUT08;
    output [65:0] RX_BYPASS_DATAOUT09;
    output [65:0] RX_BYPASS_DATAOUT10;
    output [65:0] RX_BYPASS_DATAOUT11;
    output [11:0] RX_BYPASS_ENAOUT;
    output [11:0] RX_BYPASS_IS_AVAILOUT;
    output [11:0] RX_BYPASS_IS_BADLYFRAMEDOUT;
    output [11:0] RX_BYPASS_IS_OVERFLOWOUT;
    output [11:0] RX_BYPASS_IS_SYNCEDOUT;
    output [11:0] RX_BYPASS_IS_SYNCWORDOUT;
    output [10:0] RX_CHANOUT0;
    output [10:0] RX_CHANOUT1;
    output [10:0] RX_CHANOUT2;
    output [10:0] RX_CHANOUT3;
    output [127:0] RX_DATAOUT0;
    output [127:0] RX_DATAOUT1;
    output [127:0] RX_DATAOUT2;
    output [127:0] RX_DATAOUT3;
    output RX_ENAOUT0;
    output RX_ENAOUT1;
    output RX_ENAOUT2;
    output RX_ENAOUT3;
    output RX_EOPOUT0;
    output RX_EOPOUT1;
    output RX_EOPOUT2;
    output RX_EOPOUT3;
    output RX_ERROUT0;
    output RX_ERROUT1;
    output RX_ERROUT2;
    output RX_ERROUT3;
    output [3:0] RX_MTYOUT0;
    output [3:0] RX_MTYOUT1;
    output [3:0] RX_MTYOUT2;
    output [3:0] RX_MTYOUT3;
    output RX_OVFOUT;
    output RX_SOPOUT0;
    output RX_SOPOUT1;
    output RX_SOPOUT2;
    output RX_SOPOUT3;
    output STAT_RX_ALIGNED;
    output STAT_RX_ALIGNED_ERR;
    output [11:0] STAT_RX_BAD_TYPE_ERR;
    output STAT_RX_BURSTMAX_ERR;
    output STAT_RX_BURST_ERR;
    output STAT_RX_CRC24_ERR;
    output [11:0] STAT_RX_CRC32_ERR;
    output [11:0] STAT_RX_CRC32_VALID;
    output [11:0] STAT_RX_DESCRAM_ERR;
    output [11:0] STAT_RX_DIAGWORD_INTFSTAT;
    output [11:0] STAT_RX_DIAGWORD_LANESTAT;
    output [255:0] STAT_RX_FC_STAT;
    output [11:0] STAT_RX_FRAMING_ERR;
    output STAT_RX_MEOP_ERR;
    output [11:0] STAT_RX_MF_ERR;
    output [11:0] STAT_RX_MF_LEN_ERR;
    output [11:0] STAT_RX_MF_REPEAT_ERR;
    output STAT_RX_MISALIGNED;
    output STAT_RX_MSOP_ERR;
    output [7:0] STAT_RX_MUBITS;
    output STAT_RX_MUBITS_UPDATED;
    output STAT_RX_OVERFLOW_ERR;
    output STAT_RX_RETRANS_CRC24_ERR;
    output STAT_RX_RETRANS_DISC;
    output [15:0] STAT_RX_RETRANS_LATENCY;
    output STAT_RX_RETRANS_REQ;
    output STAT_RX_RETRANS_RETRY_ERR;
    output [7:0] STAT_RX_RETRANS_SEQ;
    output STAT_RX_RETRANS_SEQ_UPDATED;
    output [2:0] STAT_RX_RETRANS_STATE;
    output [4:0] STAT_RX_RETRANS_SUBSEQ;
    output STAT_RX_RETRANS_WDOG_ERR;
    output STAT_RX_RETRANS_WRAP_ERR;
    output [11:0] STAT_RX_SYNCED;
    output [11:0] STAT_RX_SYNCED_ERR;
    output [11:0] STAT_RX_WORD_SYNC;
    output STAT_TX_BURST_ERR;
    output STAT_TX_ERRINJ_BITERR_DONE;
    output STAT_TX_OVERFLOW_ERR;
    output STAT_TX_RETRANS_BURST_ERR;
    output STAT_TX_RETRANS_BUSY;
    output STAT_TX_RETRANS_RAM_PERROUT;
    output [8:0] STAT_TX_RETRANS_RAM_RADDR;
    output STAT_TX_RETRANS_RAM_RD_B0;
    output STAT_TX_RETRANS_RAM_RD_B1;
    output STAT_TX_RETRANS_RAM_RD_B2;
    output STAT_TX_RETRANS_RAM_RD_B3;
    output [1:0] STAT_TX_RETRANS_RAM_RSEL;
    output [8:0] STAT_TX_RETRANS_RAM_WADDR;
    output [643:0] STAT_TX_RETRANS_RAM_WDATA;
    output STAT_TX_RETRANS_RAM_WE_B0;
    output STAT_TX_RETRANS_RAM_WE_B1;
    output STAT_TX_RETRANS_RAM_WE_B2;
    output STAT_TX_RETRANS_RAM_WE_B3;
    output STAT_TX_UNDERFLOW_ERR;
    output TX_OVFOUT;
    output TX_RDYOUT;
    output [63:0] TX_SERDES_DATA00;
    output [63:0] TX_SERDES_DATA01;
    output [63:0] TX_SERDES_DATA02;
    output [63:0] TX_SERDES_DATA03;
    output [63:0] TX_SERDES_DATA04;
    output [63:0] TX_SERDES_DATA05;
    output [63:0] TX_SERDES_DATA06;
    output [63:0] TX_SERDES_DATA07;
    output [63:0] TX_SERDES_DATA08;
    output [63:0] TX_SERDES_DATA09;
    output [63:0] TX_SERDES_DATA10;
    output [63:0] TX_SERDES_DATA11;
    input CORE_CLK;
    input CTL_RX_FORCE_RESYNC;
    input CTL_RX_RETRANS_ACK;
    input CTL_RX_RETRANS_ENABLE;
    input CTL_RX_RETRANS_ERRIN;
    input CTL_RX_RETRANS_FORCE_REQ;
    input CTL_RX_RETRANS_RESET;
    input CTL_RX_RETRANS_RESET_MODE;
    input CTL_TX_DIAGWORD_INTFSTAT;
    input [11:0] CTL_TX_DIAGWORD_LANESTAT;
    input CTL_TX_ENABLE;
    input CTL_TX_ERRINJ_BITERR_GO;
    input [3:0] CTL_TX_ERRINJ_BITERR_LANE;
    input [255:0] CTL_TX_FC_STAT;
    input [7:0] CTL_TX_MUBITS;
    input CTL_TX_RETRANS_ENABLE;
    input CTL_TX_RETRANS_RAM_PERRIN;
    input [643:0] CTL_TX_RETRANS_RAM_RDATA;
    input CTL_TX_RETRANS_REQ;
    input CTL_TX_RETRANS_REQ_VALID;
    input [11:0] CTL_TX_RLIM_DELTA;
    input CTL_TX_RLIM_ENABLE;
    input [7:0] CTL_TX_RLIM_INTV;
    input [11:0] CTL_TX_RLIM_MAX;
    input [9:0] DRP_ADDR;
    input DRP_CLK;
    input [15:0] DRP_DI;
    input DRP_EN;
    input DRP_WE;
    input LBUS_CLK;
    input RX_BYPASS_FORCE_REALIGNIN;
    input RX_BYPASS_RDIN;
    input RX_RESET;
    input [11:0] RX_SERDES_CLK;
    input [63:0] RX_SERDES_DATA00;
    input [63:0] RX_SERDES_DATA01;
    input [63:0] RX_SERDES_DATA02;
    input [63:0] RX_SERDES_DATA03;
    input [63:0] RX_SERDES_DATA04;
    input [63:0] RX_SERDES_DATA05;
    input [63:0] RX_SERDES_DATA06;
    input [63:0] RX_SERDES_DATA07;
    input [63:0] RX_SERDES_DATA08;
    input [63:0] RX_SERDES_DATA09;
    input [63:0] RX_SERDES_DATA10;
    input [63:0] RX_SERDES_DATA11;
    input [11:0] RX_SERDES_RESET;
    input TX_BCTLIN0;
    input TX_BCTLIN1;
    input TX_BCTLIN2;
    input TX_BCTLIN3;
    input [11:0] TX_BYPASS_CTRLIN;
    input [63:0] TX_BYPASS_DATAIN00;
    input [63:0] TX_BYPASS_DATAIN01;
    input [63:0] TX_BYPASS_DATAIN02;
    input [63:0] TX_BYPASS_DATAIN03;
    input [63:0] TX_BYPASS_DATAIN04;
    input [63:0] TX_BYPASS_DATAIN05;
    input [63:0] TX_BYPASS_DATAIN06;
    input [63:0] TX_BYPASS_DATAIN07;
    input [63:0] TX_BYPASS_DATAIN08;
    input [63:0] TX_BYPASS_DATAIN09;
    input [63:0] TX_BYPASS_DATAIN10;
    input [63:0] TX_BYPASS_DATAIN11;
    input TX_BYPASS_ENAIN;
    input [7:0] TX_BYPASS_GEARBOX_SEQIN;
    input [3:0] TX_BYPASS_MFRAMER_STATEIN;
    input [10:0] TX_CHANIN0;
    input [10:0] TX_CHANIN1;
    input [10:0] TX_CHANIN2;
    input [10:0] TX_CHANIN3;
    input [127:0] TX_DATAIN0;
    input [127:0] TX_DATAIN1;
    input [127:0] TX_DATAIN2;
    input [127:0] TX_DATAIN3;
    input TX_ENAIN0;
    input TX_ENAIN1;
    input TX_ENAIN2;
    input TX_ENAIN3;
    input TX_EOPIN0;
    input TX_EOPIN1;
    input TX_EOPIN2;
    input TX_EOPIN3;
    input TX_ERRIN0;
    input TX_ERRIN1;
    input TX_ERRIN2;
    input TX_ERRIN3;
    input [3:0] TX_MTYIN0;
    input [3:0] TX_MTYIN1;
    input [3:0] TX_MTYIN2;
    input [3:0] TX_MTYIN3;
    input TX_RESET;
    input TX_SERDES_REFCLK;
    input TX_SERDES_REFCLK_RESET;
    input TX_SOPIN0;
    input TX_SOPIN1;
    input TX_SOPIN2;
    input TX_SOPIN3;
endmodule

